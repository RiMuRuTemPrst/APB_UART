/*******************************************************************************
 *    Copyright (C) 2023 by Dolphin Technology
 *    All right reserved.
 *
 *    Copyright Notification
 *    No part may be reproduced except as authorized by written permission.
 *
 *    File Name   : dti_apb_.sv
 *    Company     : Dolphin Technology
 *    Project     : dti_apb_vip
 *    Author      : phuongnd0
 *    Module/Class: 
 *    Create Date : Sep 11th 2023
 *    Last Update : Sep 11th 2023
 *    Description : 
 ******************************************************************************
  History:

 ******************************************************************************/

typedef logic [`APB_ADDR_WIDTH-1:0] dti_apb_addr_t;
typedef logic [`APB_DATA_WIDTH-1:0] dti_apb_data_t;
typedef logic [`APB_STRB_WIDTH-1:0] dti_apb_strb_t;