/* 
 *----------------------------------------------------------------------------- 
 *     Copyright (C) 2016 by Dolphin Technology 
 *     All right reserved. 
 * 
 *     Copyright Notification 
 *     No part may be reproduced except as authorized by written permission. 
 * 
 *     Module/Class: dti_cmd_dec_ddrx 
 *     Project     : dti_gf28slpd4lp4_phy 
 *     Author      : truong 
 *     Created     : 02/01/16 16:41:01 
 *     Description : 
 * 
 *     @Last Modified by  : truong 
 *     @Last Modified time: 02-01-2016 16:41:03 
 *----------------------------------------------------------------------------- 
 */ 
typedef class dti_sysclk_seq_item; 
 
class dti_sysclk_drv extends uvm_driver #(dti_sysclk_seq_item); 
  `uvm_component_utils(dti_sysclk_drv) 
  //--------------------------------------------------------------------------- 
  //  Properties 
  //--------------------------------------------------------------------------- 
  time duration; 
 
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
U+iZuiIeD00x4HF5uOWMFCFs5DH0CAMj/dTM3IbIvzpYq/tb3F2GTw8/bL3A1toY
Lp7DOAHj47LsBB7NlwjsEPCVD1m0xgpnYQvdCJWqxrIyEYh3CFCm/YxNn+qbtDZI
AQ+hH/gc6PecfM4EyT7fFMdN9snx6YUUZxq3OyeUzw1L5a6UY88d4g==
//pragma protect end_key_block
//pragma protect digest_block
981gTvi0x0KV94KkAaUhYeuxXk4=
//pragma protect end_digest_block
//pragma protect data_block
SwKqEuiDBYo6jTqjMHedtlhvIfA0k1dtt2lQIRyeKODTPu3tzEv2LGhsfTtOknFq
dRVU6LWPQBrVm4wiK4TqTnaNHZ33r1kleairI5NQ8sdiqNDEQJ7SafEinYzgQ0H3
alCuAd2TuJEbeBQxcDClP2TNWfxmGSBJReoo7ub7hYdlx+uurHZ30C85qcTgZcxO
4I/JDYnmuscbCA6lkp72bWbccUqYKUHNIJ6VXTUYFgYeOn3OeJeqsn3p5IJXatOP
Ikwx49VekLsDSxx9ExQMXBxKXT/gDGd38Nfiz2VsUfPN06I0V73kvcmW4BxeoHAY
PdNtcMYIXrZsL/frXAIa/P9brS2xhyCiHnXJBZXUi82bm5hN2WS33YVUyiKZKvzR
cb/ZrzQ/w/vxrCq32HChPcD9I0ngGbC+PiuZeeoAmU/Q0xRs/4LC8M+9L2aCnZev
TBkjbotWQbYx798FdAkx1h7ed/2Hjo3qyrH42dnjTEeBgu0P/Zfu+0P+rt2WJ/35
OcO3O8qgKvAwNrg7AW/0gcRHDIQHVe/g5HwtHrg/vzZFACHxnPE+ha5t3H1tBmYI
Eco60sAtN6YJcTUUH26lIYZvfXA2jonberjzjffZKEgHfpujpVEsVjyylmqfW0lF
YEfGjeWAhoFp9strMOwHWNwW1sVMi5cjYOl/vASQ+6YDsyZSiHm8Ya69WGzLTgiJ
NzT6mvJwl1S8OzmHaxfZeHcwxquKDM4KdhAr5QjRdP33Fomy1CzE9G42MXm2AuGw
upeEgKA7V7/ntL7sUOyt5kCEnovl4VfEU1o3afIAChQotrS4ohfAFSL+uTLhbHhV
wjTqa9fE6tHfwtDT74K9Odd0GHNRYU0gWbEDGvJqNVUZoVOGrgq+9hiZECKqv7LN
D6QIqrFMm1VtEN3JeqkfmD8GjVG/KJNG0IDOV0nkco6g51dHY44ZmEW4a9/HzMyD
hzyr/y8mkIec2q+2es7zd6ia1P+5/koblq4BNvTUCUoUkHXji6Ly1r2EXYLP8A4J
Re5xeyLJIjVEpRNueaoGiKRoJVX5ncZnN2Pt44+o9i/Tfr0TLKmx2bwBV3f64EXK
7XAueDmbXCECPmR5l1HFprSU3UqypIAZFG/62l8M9Y4OQwikNydCEsbgJiC7OowC
RfEp7qr5GmDYJPpBX/aJXfhJUh4Nrqf2iJTL/UVUmVlcLHUTOGDTMAHokQc/JlZo
O5G9UCWtLKR0awuc5/nj7szndmTBCg5mfFFh35WuHgxMlo7fBPKMGCW7FTcF+RXh
8bXWDQeb2yZ9hUkXUwWOIvieglHqyEz7L23PI8EJ/vMecBBbLL+dtZ+7+xD6I0oa
rppRY7xvDB+JVaBvTrJuQY+nFWTdhueY/Xurs1FZoz/UPaOT1IEfFRWRaIS3BkaU
CG8dpCAzUq3e/8R2qbIJUXbaWJaLrCvqIFsFW6Vh0xLVXCQ0CihjXxbY+UYECeKw
zTxD0Lh1/n0rSKVm6+h/Ezrk2HgLYl6JO4M4uX8Pk1PHUH9/5GLa++QvOw1s3XMz
ntP+Vl2ouum/sVV3yyFbKZE6vTaFwFzUzct2huBk6GXyIq5bFuyWpuYHCSOoWm8M
802t1E+fBTvNXNabJ7/Jm5SzjLDuf8yn0i3Ds4LfUWNj/t5jjpDwpJPnC5nvsr4G
FlK0xCnLwxGn4aoJ2k2wWicxnv3v8JaCu47dWmOyDC429KcwH1mWYeqoofnfBxU+
C18npNu5sKLk7SgWh9uBnQ==
//pragma protect end_data_block
//pragma protect digest_block
49NDXxRoLUV6lJZtLI7czPWZceA=
//pragma protect end_digest_block
//pragma protect end_protected
endclass  //  dti_sysclk_drv 
