//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AMfV90nN2FWN6R0sYKMufgFgF6Cpr2LyuCC37IdX5zhSagv3ir6EnoTWqPeja++y
T6HSkt8oB5U4lNbYvLtNXCfALoO2sus5nA9LlNkJVXsNOisqOvdNvdEDHiyhfMi/
V1R/ErTPSGQRRwdCgsudcneRwNYKmX8xGwWdTFUdyPAkNOl5SXakQdbkYMgNeOAh
+jNjrUUTtj+OkaKcrLCRui89Ii1/juStsuh3kZac4Q1GsyD3Bk4UJ9K/KmUSY7+F
4g9+KZbI4Xe6eNDrDqhlTC81saiZtLrk3omkr/qznYKEgb5yoZNCwRw/v0JcYZoJ
ngBiX61PcDroXuFBNzNOOA==
//pragma protect end_key_block
//pragma protect digest_block
J7/AyNczdHu/TR9k6qDeMPJWxho=
//pragma protect end_digest_block
//pragma protect data_block
Nli+OtnvZX27Dcx6Rxk1KJFJAAvtpByx03o7GxC4Nz5MrUPcLVbHme8kCW3w/EZW
a/O8t8r+aPT+w58T9sehpKrGvI01KixnPV+bzoBZqHa+7MP3QK5QVFLsAKhwN166
0qATycsrxtGZbHj4YUGkj++E4ZxMujN3ONgAKjxplsGM+D0PBbtUAXgQiZ5Zh0z2
j00YTqcB//chiz1Fedfr6o8ohqdMjbhqPgCgxWaT0pDpVXhtCfBwmlxWWtU0+42g
X03H5qXybm0XoGF6JVQAA/JpXnNhjmd5AopebkMKgdcupZbESYRgZQMLTIFA6VHM
UY78OZMG05NUmeA72rkfKQ==
//pragma protect end_data_block
//pragma protect digest_block
mksg4pIqtVSg/1rMGZO42iCpCJ8=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
Ac/ddSUpPH9zzvMIz9A0yrL5BNkl9uv3CUkjxpzABXBWzp9JI5bgyAiFM0zoDmsL
Kqj/nUAr5uYHNMXXYOTVWjRLftePtspwvKO1Y6aDNj+FFrpJDwXHMBP6+djGZ3wA
NXSJuiomhr0HvSX3bU1rTDv2hb6HU42rMVnzQGB5OfSfwiA/kiKly9KO3YSn4qC1
u595Jpe/XHRZ48rQYIGvnFiOkbVPPD+VLkuF9HmFhQafKCgCvbLqDw262dLgPhtM
X19EAWqCH9k8SU4R70eDT79mSZqVigS0oRsBplehxv5fNi2RRDgv1I1SF1lVBaOI
P0t6YvJ+Geawd2h/6zxQYw==
//pragma protect end_key_block
//pragma protect digest_block
LCy6y3m8XhUZs7S4FZGu5N7n0Hg=
//pragma protect end_digest_block
//pragma protect data_block
MAXe2/7YQLQWxf8Cv9QLw4tlj+iJOnMQIE8v0pGH7QaQqI5+EdSVzU57GnlQA+tk
AGBLM/jFTN0rHaAr+2JV0ge5gos/eZXYxw5ZNCaqgIwwt+Crpig7CKTscLseUr6b
o7zZKmlQTWQ0ejuWNltP4N7KnH8vv5/Z7/WKb3tojI+abJ+H5A0fKbsA30RHw17f
XUJoJO5s3SHGykRbDhkMuMSzb+F6BWH5U2Szv5N+Bj1mUyWC0XTsFmpN9WLvGpIC
DL3HK5LhhK+6DwuZvOm+CGUlOJDKpFMDICorrgN6zQ1rVbrBIK1m9OUFnk/3Z5oJ
YzepA8tda6sKZhMM3w5lcA==
//pragma protect end_data_block
//pragma protect digest_block
kr5wq6IWTJGsglXt8AkYJIlEa0E=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
A08aYM7sE7vjNZ1kDvNg2RmPRKOMyqkPg+T/YnPNFuul6h2NXUdTDsaKgvdWw9K7
iU/pwEkX7KZeCUYh/F8M6IhmEPyLB+lumUKdhfa7Kjm41SQdQIMGpK2cQG4agmTB
2Cra3B/BahQw2ZLMKe3AX/mtBb7HlvUqb1+tBM/52WHV3yNplMyRjb+Hdn7pMeKM
8fFer6Yn+UPXNxAgvBHxsjEV5uSyGNtF1t2GSpkhOx74vlVgDmxAKsehNL2Fmc1U
9UN5AaYL5R6pfyrW/RIENQOk/JbkUsEUcH+cvXBuX/RcSvl3Bo1B/bPp4idt+LZM
X/YdsrWwFCu8E0FPjcPXXg==
//pragma protect end_key_block
//pragma protect digest_block
04v0UEFat3VxgWFartx6Q4wrFEk=
//pragma protect end_digest_block
//pragma protect data_block
XSfbRH73tDS/vyzsAkj0y70Hd0V22UUcKoLcJjuZlqRAxYKmgz6UBXaCs3S1qJiK
nufPoTfxCY8EwBE2BinNLvQZR2Ej3EzMJh0oIq7mxlpedQIDbIM548J4x4JAkQSP
YHix26K0XfSoxBw//zJUQ1Z1+Cy/mh/v9oBEtqCWxOY69S7dahrQvpP/qQeGZOIv
mQURPJVK8/0SdDskOLoqO0hUMyX3xD3mN2smgaTcElLC+Nwv8tRDJiDQvkR3hzGq
QpNCFiTCULEVy9HeTpm/6qodBypE1rwOZ2wCcru8dt7kQ5WgPJBJOuIc0u0rBME6
5IBnaxvB6TjP215MZBTLMw==
//pragma protect end_data_block
//pragma protect digest_block
/c3fEm3kA2lZuNP9wKJlUd9e9aY=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AExuwSfEc7mUF22h18UIHFvoH6dyvDsITonZjRaBP+GUjiudELNaFzt7701c2mfQ
seKttbIS1fjOdi1rHvDrdk0vwi7OIeOA4SCDugMAc8o/vMmTmkWZhwkCnbziSnMY
bncOmNoTniWLVEzzQI2wj/BA6HxKjHHLrvlJPbgkNZq4S59rIc1x3q5Np/FJErH4
8eisUQ7cjBuAFW/4uh7XXMK6t0chsKyKwSZz3RbKzjvmQl+jAMSOn6rnwOEUMM+S
MbXjAZ+W6Y1ncan0N0BSbWy2+q3SeGIKVteFSgHSm1O5RUASRcMSopAvC+C3Pifl
CJTQ1Un0EDYS6XnpTdyq0A==
//pragma protect end_key_block
//pragma protect digest_block
wlG/FdjLyA/GaVwkeGRCaXYXRRE=
//pragma protect end_digest_block
//pragma protect data_block
OeQFi2c0HK3T9I5BxLJdFl+gCRti5+3y++IKQ2CqxH81Ui1bjJzjwPsadoz08v0W
scyFiShuslEmK6GMOHqYLGWZpd2/aAJurmA+4JHg97UEzWFL3kHZ/lnAOZ3AqBOS
LH00eqZL3jAb9K/xG5HU9cf50a4yqr4gSbPPCesin56opKJOwpRh60+qhJrPEFC3
pKQLEhctzOCGja3UfsTq+TQdkmuWzHQIxXqwX5zONg9wKgNwIioVtdE3eMm38njB
2hXib2/NUo4+FyJcLs5ov3WKnToPtDSbFCL3RZfAPU2H2nsjN4zvUiXMV4W0fOhv
EReUC5nOFuOLGSEWc5hLiCS8u492zZIVfLkfaE+C5I2OmI6qbD3bktKamNAHVPP5
VUL6V7FJFzqqAKoG/2GTb1YirJJNJ2NfTapCLaz1/gWdXEliDIjuZoNm6uvEkzT2
xaDl/Rw3KrY7Aeq4lH0YT5XV9eE2xzztvvZNdVn0hNbJfn2VXWyAVuff2F673/Ht
h5Tkf3sZE6MlJEqx6f2BGrUYgReK0+umsIoUs3GufAhUG0w6sL/kMKNR6ROtB5pl
YSPiv4gwwCMicbr2UtnqyuMi9qNV7g0Wx6PdcvxL2Xu/wvXAwgo8P9FmLUrO/iCV
KEy6y/5GXVUUfk5FkzUTK3CTVDl4f5xfO1SfIXeggJ3CUDZ/br8l5qbM1QMg0HPm
8mZ93ZNIO+o9UR70PFP72L3IkqliwaM1QB3hJu3pe1M1rZof2iW/La54SqwVCMWw
cEFIIiFYQyspENqZQaaZ4LDXcpZFdcEtdp90WgKykBVM7tF27f9Tcbi2p/yQTIwX
zrNqEJt4k+vZUUPAwRxi7cq3acCzJM71F99xORpbwjQ5ZopX1nnNTNajjOMFYVVm
gK0tYCRNJrOjk1TFVFFF3lWMGVaaFsCLpb61sb00g6xS8g+fGM1sPWTYoHzrK6JD
Rc1uERqNK9v56bAw/vJFgn7/wQUG2v9jgAUm5q98EYySDkBDpSkJ9rOOkQpzPdgx
trTuygM3eJ2ssjoM6kiR6S1wsoQo/nE7cX2AcvF2IGqKUnGxcIH05p1eaIxOfY71
rwxlZISEQANQ1EtdE6zM2fvJ00ScxZ24j0XWaYhwmrL6Ufd0YfeYxEefQTKXL6jY
ocgL2FFrsak76wQgCPK8qNpaDZ0vuHcwc/o/NaAxW6ymiIKovTpZwFtOglqWAH9i
KkYuGmi7Ay+07IznlWhYyskDU8afIdmAlZPpZDnndrpNBkeDBX2owPFxa/OgsF3a
ylfsOvnPjbpwaCphiCxD1XdfwSNMYOi20G7jcZghrTBZUtO0FFOlc3a7E3tzjLze
QOlqbDLC7jHUheumaEvBFSnKJRsdH/68c24DPnsOPrK+Ri+8tSk5hJQhsn6IKEik
Qd8R8P+eaLHpIqZNQu/4N5hXYodUHKQyY/njouOemLd5PcCgk37gEgU+WpNGXvyA
LpFKVetPCyTCUpT3jr73iV7Rj+G2qYueuBvF/NyNXVBW2pONhNAKqWP6pE9jOYsW
oOIxeOgJqeQt+dUDSgF1TaHQeHsoZfXEMjlUtPermV/Ub87XEi9iq43UzgGOtx+w
uLRGNzA6EJPZoTv1IGuCLgZObNoVbw9pV1wPNRsmFyz1me1/e0XWXJX//52TIJzE
E3n5QXy0dey49HJ42aNNnM7IHsb2Q7IVhypcZnTZ7N+RCLeQKeQL+V0c4hKENlbf
QL2AUaW2W7HpkHNTRx2cGUgjGq15YoCSCPpDxTT91uXWoqCw1LrK84uRZp9iZwFs
E3MmRhasc/U53hBCbFvfx8IqZsaonZgJAQe/dGvbYYupiX6MlpI+whtQSMdsVcCJ
twtUKQg93i8J4nppoUORYCEbFUXdjr2Lkg0RcR0TUcRqTZBX0qmUdRIopLYRa4A7
f2oLBPak47OogrUkX6TiybjKj/xLFSYy0xi26p2NK+qM5sJyn1baG3x/vOk53kHm
JTI9OueeDAkRODyGTeud5Md0mn60hSxfUMr0SrTL5vT+/bCm5UAp+cUx+qBR7nIh
YvbMQkaglnQS1lBAIVVxeyDsF//nPVYaMKfbF+mrY+AtuqF5g4PErECiSqwHcopk
eZ/kypJBTr6ozoHI/u+XUpAd2eBEgAZeKiokJey0cvIMQlkh4rGTwdaeSktOchu9
zM6VXaAF3oO5c+QBsi1mQQJduH9kvWJwTvm48jwiYfL0IqTvzgNPMUO5drLKaykS
jubCiDH9SQiHWt/KzJuHUjFbA3QIR2s9Njw/uFkAiUNVFdoi4d5zB1z23QilmUXS
r9zoAoweyriVMWgfR+Cl5K346Z4CA0yqm2anZEN7jC3MCxa79Gi8hwLrrCRnRhhq
jCePvduE4UYhLJI7s8xU0Ne41x+sHHP3sXiXMxuVv8SP2qq9HqcUNRXRkFu8ZycL
BWo4p23hD4iQI84PYNvs7fXfVO8XihHHfRaZJQ3uSIio4lN4rsRF7VGcEJGvlkcQ
H9IPKBWsnvDogfT97oHzGGtN2x7pgJlHbVc9AWJ/hqFvMT7Om9/aYP7sU69rmtHK
hjyOSe6CEetNcnp4YCUMDT4x2vPsT2KtC1WuSxraerg4S6SMEJUP32qlB2FU23sI
r8+trE63HywSn8NGwcJeNpiWNCOBE+RFBSM9VExjihPHjr9Jjq5pLPpOSGNifep3
IOjJ95140eU+Jj7lERhzPdMdDOpi0igBx8ZCyyZYNPaiWVNbSOApLiYE1jn0K00h
xSIt2FDPJZeA85q16wlQIchwUKUSND4ZPBk1PxLjPHT8SNWzHVSIDkOa/K6/8JsS
kV6X0V7yrUBpGWhXUrGxL9sUGYHU0XhsmgDg7hAUOTvRNDCXmlXDaSB13LSFZ58v
Ix5ftjeYSFM8GSYKJY7rEDD4f8E585OXZ6I/L3eqiitwOIqUiFa6e4U1zaVrjwqg
At8zMkKClu3xxlak01L7jk08soNZEDvOWiDx6bERAuW9tO1SghjNfXCSOL6HeDH2
KTKRRON9Qh/5bWmfww3ljvHGl/UlaP0iREOrTl12DUTzLf458MqwIQMqEUEQIUX1
bu2r65+YnFGewtkwkG+y8lRvYrJ4qp4/Rv8dfEcII1ho0kUPuh+rRFTSmCW33d4W
BOah4f+I3d3IVvBWzMxnSkwjqr1m6XcigQqyvFjJVh9Xxzt5WPU7i/uZ/P3kuXYQ
W/KwEh5aYzAQLLPSCIdODNnwflmz55/FWI4sP7db7wnK26man8kkQjOVBn3RII1W
Lpwjn50tn59Rx6sQ0iryDcOutw2MmKdZGleRIfdRwdLKql5LEOFKxel4LWjxMnzi
3vdFZg+JPykK0yql5npoeCnse3r/anoiUma63PQdUkcB3MHpT95c6D4aHtmqH0kT
AwSNtW5WuFITrrSYl4r9t+DfGV7YkYPDPlg/GoZ2Xf6Du5T13a66Xziszxrfq9IR
CzPHFX0CDflvK/1BCwpQpLlhD9kZPCdL9sjSUshnZr/dHlqFptvvF2rGO9JfpswI
srte9Wq2yQUSe1vsIqpcdvyNozOEvdzFxrnpkXtySI0rqnB3AVY/Gzwpuul7TlSC
xWlSLQ6Vg9r5YpZxkWkeeYrdZoZnaZH0XIoI/1OZeeB7GdjZirDXRs9kb1pkrPUE
OICClb5TySK9DtnxA/7KShBmfKt7uL7GX6zv+DHnKRbdlRr903dNgHzdTRbvOV3u
5FZgowKZygbpZHKtaNb188o42UuDyN+naV7DqaPaVjKV+j6F4gIzMTzlQjs2KJ0q
NmtvLnwtJo8m3nUmkSnsOU8LiFyufenZ/uQ6mhy3ZT2IvJu+U1xhytPPjdQaRTO/
U722aa+VJ0q/arXJLyhny3as6wJ4555ZueunnasEcolM0TlCz4o/z9X8N4wpZL+g
YUqRZQjk6ya5qwVDclEv3V5XTgiArcWOY9JvcxhBu1aJQEjLy8fdxIMebyfBBD0K
sKGqRg2b0VL5iIf9RkmsIMhYCCSJbWJBd4ObGCBnuNhPON8Eat3VVV5qv5wBKYOU
WYen4NckvMHigEhVsurbVNmSrOqx6PeJ6VlSRqWx1eaqaGZrOoOuXeqQwgOW5jv3
Z2AyegrPx3hQ4/x3F+0eZz3Yle8HkkityGrdqs1V6uAvYW9S6oL3+qp+GEKfkt6t
mbYSSH60UMQHCyeyZi5pi5H8S7EXl9fuuGtNsLHLgXDwNbT4kOG2Rd6Zjkc9LbFR
1j+BuFfEJlxWJOMu+sn2zAvN7EJ+zmTuD9h/rs0YDywWQJppOS3SlMlK7pq/lSfI
suEnDdawh4a7/OEzQF5Gjz50E3ruPqdZGjon1z0Y26aJiT7Iicc95VUgtvzTAwem
F7TBizpRuJm0EVX0c2/3grovOQuJkU5BaIOTTXJG5QPh7NIWjVXjB1d5ZhpKWI1M
DSh1wW0W1AkCwtMdXJAbXqNngVzikO9jjbVOLEG+/AHvh0zvXzSBwi5jMp2JFnNi
OahcbyBWQ8Yl+D7u9HRJHeitqYF0vKoyHJtCABMYp2HpykhTzvSEmv2yc6fxiiMW
a8xL9jy5Z2LtwIlPi2RU+Zva9bOwula+MNVPYFWISmV6J03avxBBys0PVcGv2yHT
2L9b76cNJ5AnUrBLgoxgeggc55wXMbjuT27gpGJE4kyfUJr3k1V6G41Nl3YmXT64
1AUPluH76CA+tikSkRqDws/2UvXqTuyqFJoswVv0MZkaCNtgnp10c8i8r3nEupri
SksQtCwTJALB5kV5eE5eyeGxyUPzZWf6UmtL7fN2tnDknCNdUVt61n9b36v48WSM
Gc13uMEMM39Ga9rad+E4MSS17hy5bIkctTNjZtCezDD17WooZUy8lysfcXdejA+E
kuGr5kcCc3N++jMkTtFRv32zczghDzIdL32X8AxpEUx8QlNJIO1aaQuy8qSufGFL
7Zg66ZvNL8gGdNapxCp5NIWXq+y6RNlMIHJI+N2ZIyn8rOtk6/PCG6CdTZEsooo3
tSBw2z8AzX2v/FblcaiufqIiMJ+ds5S9Frty6f1r3oaSeMWKV1MG9WEZcaqnm64x
pGfEV7jlMN8lKXSbiQ5bDcoyBdb5jS1581X1yyO1JPBxXj4yPL+ba0Mv+wFt3wfA
b/PguRQuKinBGB9hx8WBb8h/A0CZHcajG7/TcWsQoGAdm0B1wdjhE+E1E5w9jtxf
r1Sl0Mug51NMC9rUCnfouG9cwmAcsBdJrBpiPB5Zb/axvxJrghoJUxO129jB2yse
wIL9dGjsDjBd0zmB5PR11ehBHyoiQ02lukxEmZLqlzN3qhNW2ykLNePXHuP9fZhH
z/87jcFfNrxeSIQMib1po47PjMLzAyOBYrPAFS7cMlzr0Q7oBnY8glCN1kUNqlB7
CLqN6PhVO/MThKI5cwQ+D8YNjc7A0HXyaAl5qlhER1TJjGL4Ww2PMIkHTFy4fJpk
giqcVIHN3nNtcf7sh0UA256K4wCf4vjuIBCOucBoFaWr7cEcqoOD64foI1f+HcAd
mrqlg47kj1rzrwrA6C6LLNn7Vtu8ybw27ycSoC3q//hkIO+CubcVBa1VNY+QDs9B
ERn1mNrb8Ne9aLhYAg4mgtnVHW+PQWmII7WCjw0juU2hm7NXs6ILb3u/KiRuu/lM
WQafl3aq0DwWc5jhf99euHNjfxBxOrfqLOATkmh/OsYV8abfHDF3JbA17xwAvUNZ
912IlVcuKrOvaRAJiUMcJAfIdiix76DC2F2Ihlqh44+5SWiA0mEFpEPFyD74KxB/
ro3LaO/4nJT5qOlI4a/+d+fdtJnlRvu2eMtMx+7Y3vmbitHx9wmBMCX0mb8PAjFj
IMCDcyfcRAkswwo5K3/34P4xer0hUs3zv0aYv4QJSrf0S1X61kaNJcU7z4iln30D
4NhXw3UebHPp08w0KfqmyZGlMU2gDkg1Btsu37UsA5kUgBQIKNffgAz60FVBx1PB
6jh95IGMJEAdvoLvz/H/7GkhHyQE3Fj9F7zR0fCZ8GD5DiuNcX6mKPR7Na7djTVh
nTH9YRH3MzKffb5vsviPZzhNwzKqDWtdq99cq4vRCVHRlPDbAoxaWL4cB5jPJbqI
I+uAe0omXE/qiLsXgQMGCUuW6CxRBxMLv+8AfFJNWysmfiErXcgx6vYNBTyw1IVS
N5Bqb07Liy9DL9DMI5OA2va48bq51UbNVa1julCyLPQUa010WsCIXe8YkHzRPOo9
7i56mSSs8IjcV7gpqWrYKL5Jk8chSqObBhbnRYWRKqCBRFGOdTGO/QqgUTYLLWAK
1eGEYHBaD+X2fh8iIQPRrUBSRD7ffacydahnbWsMJkKuYf6+Oabd37tgiPxlrmiT
n0xxzWII8fSfrtYCnxuy/W7HRJq8cqr3l27lfxyMxICX9DIhlUU4RpTMUa8QhHGL
7pBPX8FCPlPUNOc3a+ImLKwDKh1DGB4KDdo/ZZoZLU5BYgrYGUbQnKvyylTATLhd
ZHdAvL4Z39QpeG5S0yaYmdWVPaSdUQPZmSKD3SC842sFDRHFo3SprXdxnRNWlzpF
0ScWOA/R3sWStBBeePBXyMdr+yk0t5aUQmp3o/lCuhMxN85fCVYmj4/tuMuHHxoz
XYRNQngToivhe22rTivEuxNrKDAf1ZbIbKmyhP5hZqdxKKBsbARIfVUVebOQ3RLr
Ubka0oG3FSXDHO8twJz3ic1Z9lGOvmCe/p2xYAu05IE6j3iGFIz+rNpiDezJWpXG
wsEy92hWqNF4Mb0rFSUOcuP01PsksFIRPF6cjBAlEM3VzBHYSF6ZFj5Y0Gw1SUoe
ipvQ1bfShQGCwAsIZjy6gvqQtaUUu0UfPuciPfu++h3pk9WK/MC9HgXPyOd4ogV0
xTj1pIzjL01165kORzfNyBEe/ONIpolf4L3+B1Pr4V5E0faK1ZBj2FESFn6apmK+
S8cgVjH6QOrlnar8C0OwYqr6b+ZMD2XsCxBEBM30qi9m87kdK9jnxvFwT1Skjfps
9gBPwjoJFmKxdGniCHdVCQHQk+kRpT+9rQYJHlNjBnNwHYykGEmOZTUV8GOiYYz9
Qkz7A2vLWmqbHZdmKRgwkQJcGjkTELQmJXyiPM99H0dX1q8dvKLfhyBm6+tsk/FW
XCsx9tAD9gH55+xliNI5H+dH2nkRVTt1eHWI7x4TXDWjCs03yNi+GGHgh+ApG+fE
lrDraggFhpyD3K6oHsPcN6gNGgs0nzesRJPQAq8TrYpIN7iGEh7POb2HXbtYU5Ua
j+3DleL3f7QOwzObRFdMJ1YkVjI8xX3HBGt+T1CrdIeVGDcalAAeRdzrpbL1qKwg
d45le6Q1WLPl43dOPnm49FvKzudvJF1fcQv63QI3YlnK6KvENRDLuinrGo6M9oeT
DioPx6u+UDaUjHDngGYZyFyURpzTVQ0Kt+zBvD3VSJcSF8yrjUIY6S0gU1ttFINl
U1xpDLKEeyQMJKq6VqBlA3d7WxcSQ+4OHPOKAYyD7hHV1UF3gpmTRc2z/9IFiS7V
IGXKjPBOyYy7nhHxXxE2fr3/GkUN5W0kNw+HY0qJfnpZmp9vUh2vNxIveQ4hP2FB
The7xYnUyL8atgDSgg/gUqTC2b+sQP4lTkPpSq/ti4B3mlqSyOCKX6DdQs48U/fg
DiKYgU2N6p3u/cnE6B0Mkg5c4BFoD7xWD8+/70eRhXPW9BI0T5+VJdNMOK847qUp
Ere+VZG7E2TyBhAKazTv1ItYw14TvHWXymsDUF12xpGHR9CTOwkGelXWLiKG3yV+
GhbV7v+22o6W7Fax4YyeuxSwrmrFVfM4wigulwdXRJjDmoAckEmsththuV1T2wIG
SChhWkmkPt8mNWe6YCOzo1z41htmdEVSeIGiBD2EvwPPSZcWoF762SKZRnT5U3GG
WV7gkaHy8YbK7Q7wp0IMhJ/ot7SLm4YciEveCnvn6oUHGZ6cdL2n2likslfDQB8E
iOaRnrliT046LRcTjcrUGpNA1pPFoibUhpkv5JwWR1nSHSSg5vOy65B+5cEjOVkM
Yb6MPCvfQOJY3LGgnpWuF/aFITFKyu/JS1v52E+7jwnB28WFEtgyqFGaJtn/Fx2l
3SXkZ0KKrMYZevaIVOy9OKO9MOJpol5UfJRZoSjaaj8iW4J7nEdo7JrkMQW4Wlzs
qGYxrMUuKRIpMNRASAL5MvYHaET6lNFzwN8M3EpxQC488yOj5QYBpSrKQcBVxzx0
9AtKQM4N257lkW8hY2FSWBQZLwAFCwMnoEcPhYop0gOA05JsQsUNfnjQLOL6b7OR
UhhoQg+z/HGbT4m0+OkMwVXncTsJ4sU9dC8Hp3UVBn3ROTlS750DAoIzFUHytbAx
rbWQLFHF9tlnp/B2y38LvsoBpB3U4DEqYqVwuMdBg/jZl7sZZLIDQTbkyNJeoAXw
6lgWoG0LMtlGTMbu7u0wfgTbyZj1zZqoo/kNOmr+Y9QHYUAzLYxG+P4h6Wj0EnAG
7Bi28yqFaNvjwwMHFqSgcEz7aEmBVfUViw+KSl/sjI+qFCx3jyLUFjcFevoLkcUh
W5Hndgl1MRuD655U+iRmy9cVwG5lZTmSJ52szg6xEOUnCs60mhMOFbowZ17NpZdp
75zBB5H+5VE5FFHeGhEvlVr0rNUX/SXUeEmR8kLT+Ya7xXDMyOHAcERgsAVPvfLj
1Ml3jqqFesONojjlF8tlWDcrfROiZACqLQoEg3YtGQQ7k1UfGnnarL6QjNvXrIeH
bVw6S8rYh81DKBPns/YiGhQ9s7RBka8oFZGvzSaLb9tO7R+5QjYmbyDTInUwFMtP
Yf+h1veLwplujSjfg4Ak43Fs3rRJDkdSmVJrPD/0rr6nFX6eqrbVJUqjKAahQkJd
xsHo0W94EXd1P84bQ5COx4H8Fw0zNL60T88shZvqZ1HnG0x9FJAIi1WVtfR9UkMM
5DEi8IW1o12oGu9qArRXt7A9nSdYKXDCDMcewoPMNCqF2dM1H0MfvrqlHTCaPAE6
hA4eHfcLm0IliP1kP4N+vKEIxqXxrPRA7x5F/UKdINPqG5Gb2Jn+sXgPDWpWL20P
UibIZ/G8xGnkCVQgYM9W1KlrCRIZt05es/xGvD5dldrLUIZSVQ5NcRj42MlWeAl/
nvLvXxPN0uFAQJ1KqhSjaoy2VF2hybtimD4UgTgNtikFxKhmFvvdFztBmJvQuPQA
7CeFD3U9PsQZbIN+Om0t77kl1Jc5vUwF1rLMJ78pN5zdPW7wic+DMIWfOMfEuCC8
yK/jnzk9UG4rE+VwoOoxrunF5SVQJPDUivxUxKtb9xIqPgHLTRh8w0RnSVzKhaAn
1Npvs5LLSbDz6nk8jNdPReCXtff8cVn1cX38GnGwECKwCTY0Y6jKuUuFeegW33Ek
nSUMhwWKRypt89Z9Q1X3E1NbjIOZ5w0TklB1qIWyZd2dnjal/DvpZCwETX4+5rJ3
Tw5bRxZQ/Qzwh6/VwZHru6oXHXwggPUJIhcJc90SkX3LWelJXCLEMIFkjapA63Uw
XgDmyEUrWv/QX4apTW+VT83fpK1ISfmqpM18gnhtmlR98pEQMM1XErCf04ml8cx8
aforA5SP0FBhHHmobzqVEBtQoLpqsAWifvVt4L+9mfgR7uQVtlnEfN4XnL2Lex8h
aNrDolbhTxB1LHd0UPJEnASkNi+4QRzDr/HJrh7z4q1MQIKXECtrNCneHI8T5nrU
B1BJ6vkZyrxpiVr2FteldDJ6s4wY2jyXQhhTXycoJDHk6ghsAww95YTOvmyCX059
xYqvOGuCYoO9Kh+TC5kHJZ7W+KAhRpi02PfZB+Q4voXoqYFH6ND6LJd1apn6x2Pn
CtKwEfxM2PLsDwvoZLX8jXIfKFNquzaVKaRfx1fSSAj8FGBNLULeGPnBT8NAVVhL
Lpc44vDvn8CqrGRK6Vv4HH1D+PU2QtBPnFgYEGiAi9ROdTDt2sIUIeQsBQDIV1OI
SwmjEODuzqmIIPvlGux4xcE/Yqli94FZ21jhfY6bbgGxpo2G9jKmxC1jS07o9zUZ
IP/5DUcayIMYKSbLlZxWcspWvyPoF+f5nBVqivOPON/3wWOrsoEi8N79FQsv+qXV
4bp6rT6uHUUcVlxwCjcJUupXF0dftNJzrBBE9vNJ9N0ayQapZ8rMEdUSCt9p/TbL
ZZtaBgKXYkvdYbFgVFprc0kXNxVHrFfpoW0DvUKtziP52buCeugi3uWthe5SZZnR
EkpmozYP6UgdlePd9ZJBEo4dlbnarbdytxdPE9JRwzC3dqiuwjwlbs3mUpIRR9wi
4rw/6k3jLMHtjA+3LGpeY+w10OB5/Abxrr2kjCkgb4nQRywZDijFhFT/3346f8nK
Gzl4KcRtZvD617JKXBimLN/esG/xGAAItzsT/SfvxviFKY3EJpraUUzGbaZFefAq
orr2vlQ9yoAlH4VsY1//0IZ7PAkebhpwKSGuskBtOmh5NSPpsKAJdwZaRZBQB6Wj
Ui1Z8Kd4D71zvNu4Xz5Vlbw6/PjuBWi/qbKG27NrG7R/OQFAPDo4tGJHAjs3WiE7
izpq9Z3Jeg5lOmRT22hS7CLeGOD5UoxKiGhGeOmNL+lJGUkjyfgAWzFGSjWirxpU
lOfS4TeGOnfVhFV7ZlMTqnqryktru0jXcCRhBjdjY8NkyHX4EnMVIib/huCYuuU0
GATm0g3brj57my/dIoA2H8QsWLUi6IVW6FZXOZAHZRqw1mWW1X850nrl74GeSijx
t4tLbI84TP5BLWF9vXhh9vxOlWF+NsYNYZ67osusrJluMdYkTIe3ex238jxGev1n
oBDqQgr/CsNw5sIeqKoeWbSKqsBG9CSBnLoNA01SDZCWHjHaFmC6SzDYpuEjrfgP
Z9re4CpHf2MPs8UBWnerz/BKQpmnFoQzgbfu1r+xUsv5hLFHFBlgQHkSARurbkko
8DzIXl6RwoLWBgpch9lEzCg99G7080MI2RJOrURB1/d401sQW5JKOZkX1ivLlwBx
/CcPVpru8VN4hWOuMWH+P+MhqpqzRrkOh2bmBe97UEqp5UN6QhZ/867fxXHAKM8x
VEl6Oj2d/UkJ+Q5CCZObf6viCC3eDERllctXfpveNuPlaUMUNiUxcq5tc+utCUhP
TDPllVjPGSDdVWmjcLioiot0GJyRFeasVTtMIx8NlcUxQ9FRYP2H/OA8VuArlosG
gtAQYYsRvK4p9XoZkVYufAjmhAHRbLPkfhFJMD3lXrpznixSmUSIHt0V43tYSMxd
vAP33xvpMjh53ePzEWGEWgIsTum0D3SLEUIAeQ03WkTvFjYptWUVI6uZJCiO1cd6
ZD4V4CsYC3sYg24qm7e43TPFY+7kJ6XWJiyKHnN6Pg3uOcxHHgExAhp2fFVNX61+
no+UqFcAU/ze9CBmOjAuZ/8kMF5DWphCNruCq2gU5/m56a2SV2/phKtdKnGuP90q
n2qkwJFcc4r8sabWo0QJX/brza4Hg/n20zewvG8LRZKs5+QB+iK87TZ7jYsiTsaD
JpJozHnDgC6jA8aYnoYB9Y1sdZ44/VZ54OzIZV5+xCN/+t51zt4pokGeW0gWVUGK
rbxg8mzYBqGA+AE+lTOFLIuXvVohbUm3n0ExO/krXN/e5f+BITvwTIHMv0BtdqhQ
tLhyYhHz67H1WqmheritG9oDBm6HU8h6kux12gobNoN2gT8fquj6BhCSvkym8UcS
yA4ef/2SAF8plV+zLAwtX/9LL2FjRN1SqLKqSmjbhT/gejPd8kzARTa7wOmOAUjf
iyPMclPXwCfFBYwXayOpu8CdiHmQj/CkGmsmGCjjUYCHA9Led29s8S9yQDJp81Wn
SC97beUEvkNOMuelHdtMp3XtZKI2MSHX7HSnBh9hcbbsN/qTkvl+/RQ1PyedP1cy
bXEoJChXagpTywcYjtyexZjaIgn6vxwJDbbDvAvDLekC/yblQy0PnTHk0zvdne1h
dWnVUVAvO/DR8aHqNJWCNNL+mcR5fefr9YHhCY1fGYpzjwWZAGQ4L9+55QzdMlzX
/wsHLLAsAAPf1TwFvtPi4e0vN0wzlDMHIq8j8xIYPYqDeMVjeththnljtLkduAxs
8kvJ3TuLRThPz8EVTWyqcVzT+EfZ6092PJmgvG6QkiKT8AIhfFSZifDFRfa7FNm+
FKjGkR9L+zvyX0WNkph9F26vX6mn+DawSsRU3CNehmrmPoW9oG/MQgsmSGIN3YrP
pOeuf8dpRunJdV4R0e5Q0HdYLs7iQD4xArSgzET6BKSt1Wy1lKQQM5RPoa61XFbc
1kWU8svhc6SCMKWKtfZX1kSj/djQgJOUAI2fRyF0/ROb3CKTMGsKpwgsrjNe/Blb
HzmHk+A3fj6eQpSjhSGWGm3wZlpv2axs4Qg64nw+RZoH+C+ZH5wJlNRlbJAo61r0
p+CaAKz9FnS/isMQ3R4r3UC7CEvAIsyLtedZdpubytPAeypP1RQ0crlc678PJefA
RAyvFsiM70Kcm/lAdLpCznmLo/7Z8ygBU4CL/qfCjnRcTj/tRlZledHlvTyJTvjf
3qFfEjy7pPbtaaivs9791eBXwCx7seRfJ8bXniPsIaNYkf2sCFPa62mbs9sqoSEk
euKDocLRSDCuHV3tAFQJfNxFERLfI1j/VVuOn149IAwwMO6YsTxIzLRmgcMaC08y
70nrX35JUWi5vfTH/D0iBlVFAbOm9KrFIYrkhqMQYJmqoatJ7jZWLbRYEUPSgWYJ
3eSOeiRK7RhmgA/bgZXV2BrsfMtMWOta7+LM0B48qlot0zeNm4ndA0mga6hcFZQF
VYLpBNcdH6EtY3AXlT75qnFsR4B8/k9cexfLU5/lzaMogDDJVU7jGbx4SZjE5FO8
TilrtYp8w6cv+Txp5gPMyqYcQ3JyZaCuz/LYGlgsQJutS9z9c1+P+v64o/IHdRFM
wJlPgLeY7hpafBJV0qbUBXo2zPW3AmIWyNCyEjMLLL9heZudvZ+OKbzHPqqvg+Pn
lhdZsB0uL/O7uwrb+1gU9zVtCjtBCnJd4CrsI8GWXp6eaBWZwtSuKZ6KKKOTQmyH
yKkzZ61CGgOhmJkgeH1qnm4l+xoGyDq31YvZrjju8NauO54UZCNYmXpyHWuihuz8
vTfffkIVod8UrT1q+DYqZSKIdSL1pSaDNugbNlMnoVqDhEpWARfY6KJWsBXJtSMc
MGXVhoOxf4S4kgIgCJ0o49kRl3jBLZ7Z0uH2J66TBAdGdzDuELDWp3BDoGf/lvWs
o+pDZu/Z0Chjbk72acVU1v8ZJw/V4mWxm0L1DEltCPSJ8QLWgnwEcC5dsqQ5bBLH
6LJSnZzmp+VYIu2QY88+X19vSfdYr5LRoudw1N9y41WKckA8+E2WtegREuLTd0c5
UGsqVDA5v2+lgsVtNJzkMmelhFzNyQPJzUahfTmGpN9Pr0+ox7rzWjPLb4EFn0a1
cEfwJB0uS3ylVpsCqegZ1nH6SbKlCCqsqS53sKGaHCVQloGdwXYqbLKYMoKj4gtL
19A+CgN2Xu00s6KztH4kpmWz/3sOvmIOAdCMbsym5WYTdgYXgnh9v0Q9TZEQUgGA
zTo2pHkW+gp105SFtau5kW5DKhm88+j/D29qXqr0bP8AA+I20oLzTKJr5o3lMTyC
YGQXngAEzKQrd2uo87qPWkD431cgzxtMbgFBaN4XZvOOYjPh52XZj8hparYP/Lhu
o8RqZfS1kQZmOsWTTOlEeiF7QmT27eBARxughoL/HI2Jzj5H9W4B93VbOzBzqpX7
F7Pn7zRfhSBKzKeuUwvLixmGaCWifQ/3/tjDbNpx5mCt9jK7chOQn41qXhnu5KOK
LcbzgZaaTi2PUCGN9sitk+hJ2GCQshs2pQCVJj0hpy2SHUAh1hGQVdb8/Yd8jC02
4CJrtjuBM7LkhWpbzxPzr+6RXm3PbUEIAeCGaQOjDo+3t0vX57kXK+k3Qzuks0kf
/xtn+sLpFUnJ/J0NaJ6xIpRmoBiRM3OsiIWdCs1m+43ZZj/Q/zWIjRnx7eSVsUsv
hObQnEN8wOAeI1YOGGWvGaJMxpbwyNX+lFloWX60YmYgDO2VhIO7Kisu9AlQWUpK
bPsNx9eTIdIP3oG6BJOi1+TqJBfHaMioBnfpTTuYShU2FEgBtFXiFCGE/2/rCnUr
Q7k9teo2CrbIOCvofm8nbMf2E0zA2FkHxCJbjYKSgEYF7k8yh8YR+wCjQz0+9PKG
3wCV8UWwvtHcdr0u8ctLFTlWZRPIXE8cbSYmDKN6LGeWOMkBkHntvHxujnQ/izCf
qbE4Ib/tMj44EPK7m+pa7G80N9WD/ZnhmepP5ESrFjAZLFCrk8qhEuet/EXSJ32Y
OnuQqpGR4w6AvvbpSkR5/+DhYUXGIC6MOnRoqboXN+HyRcnKpARfyTWEY9cI52uz
a21wvXGcVVFaGpk+5U/ucPn7+N6hsMEHnoSCfcvZk/pLfrJc4EhabOFRNe2Y9OAk
zkaEonXncrOkoaqphm2WFfFJ7A/Vx+qO90aliAmbUEfyJ+MrgHtkJWAmNLuW/LVz
kgFzVa5xCXzYJIIjCc00cTh+ERtWYfpf3heUv8CCdpDxScNFuxtbyX3p1cL8lN6z
sSV99aDdToIqMaMe6i/j2GUyYTkNgmbhtus+6tlpkDisUpFpyaf9VKZCDXeGY7vX
pfynmpK5ILNRj038aiXn3CgY2IQNRnXFyzV/pkN36YHCjtILFJE9Yc15I6+lmAgn
9l5yqMgY4zGRC2Ve0/Ql5GFs6NscNVtaY8Hb4eYAqlwJymhH/lOqx+5VV7uvzXi0
zc5qovlheMZrfEHpQpIPWj++ebSFbgsKDTQj8GPOIuWcTrH00o+NWiyHiqz2Ajxw
Ys2U98DXf8ve/2NMd7yj6tJMK8bnGZAsQmm5RtQDyYKuOJhIMh4InWCbWRtnwMI6
R1a8YMIhHRFIn6ix8Q5jPF8cp9uLqEBJaSqT3ZG+VwfgW+nM3LhfzuPqhuDlvunQ
U7ffPhrN7IvCFPutfhSN7f1AFiqg904jpioeUT9mFDKR3zHGyPu5qPYn2SemT/8r
kbsw6Zbuto9TuQQd2QK9CcnEiSKO/4x7+4duaoZK8NmZpuQl7IPAvCW0oCCCInAu
+8TvsCo+ab0PtSoNZa/UEHyIBpaadQmIvD6b7TxDuTRy1MOM/P0RGlR1VDhWXyLy
Yhy+ZBzIQDqxi5FoKWPcRT7joUE4DPWTPA3Ygh9LOkjn5YeMFvG6McxmCjg3QTsP
D1lvfjhBq6JjMJr96l4Bd01cOes9r/XXdKxqcd28RrHf4ITmgA1trF2A/26f85Pn
zy1CEtY3ZRA2M0iw2ibb75XkysM1IXdSlPBH9Qgnwx0OxJEMNNUn0zMoMAA7zA8P
eWtMpE6/Zps8O6CoAzPpDLhurjTXaXP/f5sRviOADpe+/hrxvjaQXaL+nU5lJdvj
xZmHcR0FRsh2cfh+/VUT3hYY/CVreXkOYvrJ8YxRZUf2BHafeP8CGskuuPcV4Aun
JFAvekZA17gt6z0UjsDPOBWRwdM+8BZve4D6XMwtQmwksplCPIT6Nmu0jQdfmXo8
gOL0JIXWY0S9KBMaUElQ0cV//yAlEobxyDAMcrmADmHsUSUPMmOp41TxEOTRCMnz
rY5ZTkGlVGjO+8EuHnZumPyJr2OG1fSpHcGdo+dv/ujHKk3wqqeVO5i8TS8wH6UW
cal+ngI0b2WxO/lay4rN0w4oIeg9Qah9bgL5HsGdQKkdM+iiRk+ICCDUH4xaNTLw
l7e4y3c3bKic3kZVgybrqY1//fwnnAp/+8VBDoUft/TynTt2uGFvoY+ZfpZJs3CE
TdfBomcmGKqish/Oar0QzbLuomnS+IYlXmAv6rc3nbESDzc4LIauUyKbM3W0c/Xp
cGmUNPV1XYvU/KOKqByKNhy483sIcXLBJ61ghHRDIOA=
//pragma protect end_data_block
//pragma protect digest_block
0e1CVJ+4b3ZjYPhxhSyS7MtWNsE=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AOyTt0N/K1ua3Tc3L7L80981oIwhjhLJVR6QLRAyhPWVO3vnmnpjPRrqMQ8knXQN
ylam/LdFdu5vjcyZVensUZHG8GtVuxVenRW0ZhxmMOszG34a4lCgaS0BnIiKtL8z
yFuD940jqULic4c5u5GSq0wx9bN6edL8Xvd4AgRRxLMZxyyZtFRD4W+i4ufkTo6C
E5HMtaIadFvSHI9JLAUKpB2MxxKLuLT7IBDzWCUVt4w+Z7oUpBfmSi2BUe+Gurqc
VereBBxpgqc2Kti38jmN3inpd/kHH59uWi4JW0ejN+hmmgW5g6AyD1xvWGfgfhVm
G50sdYyZHdeyA2mOVV12Bw==
//pragma protect end_key_block
//pragma protect digest_block
XdVGduk+Q+zbqNJz/9/D3oTHNeo=
//pragma protect end_digest_block
//pragma protect data_block
mBVVCW54nS8KKDruKajYi9DzObva7VydepuKJP3hYOx/k3GyeBM/EbD0dbz9O83v
C1D6QuezJ0cX+SZWEo5J54SSU/dD58KQRnOwn43kVCtb2Ic0BaVjBZJL/lts9MeC
t9TZPD54HKXH0UUCROxLh1kCXAj02QfheeZSBp01zbOWfbXyYtFbaZHmw0Ct342e
3ZmkSMoaB1QaeYZHNpKTUKiZSKSr3MOiqQYSCjGKTNIFpg6tn8Q+CL8xgGpH1e19
DHqlkGtkV7kVYkXwoAoSN0TzGezu/ty/O+BgLEzbIBUR8AJF4e76Z4IuVaFtwPEt
tXjuUVZyo8U7PVQ8VesnRQ==
//pragma protect end_data_block
//pragma protect digest_block
hyVdWBZCutQ0K7AJyea0+3zWzZ0=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AyyYsKNRRso3jUHO4HOcLVF3qQPaX8M2u81Lx0xSw6ezow7nqLT9WcmTk1+IOeJm
9P6RnYpCrYT2WomgCfNBjpv7YSzirPcIOn/7877sKzDqUJxzaDhiHdTImg3yjTro
F3IRBqSJpd33uFIlDgcVHQ/ZgtJjlWh1p7DdiB05YGfObtoxznjHQFxjZrfuq01g
DjH40Ey6FsrOX7hiOsISOLX0tWW1sqiU7VD6SebhQNp1boFBcGE48Ekz9qGEnQRX
5SyeusTAJIGGbjVf4krQ1/uqC+lLaVTrlQ5Pw66Nl8npkvkhhWzUxerAZgDVCIkR
ykuhYInuBigaWWe26+9Evg==
//pragma protect end_key_block
//pragma protect digest_block
EnEM5Dw4qoeoqcPCLf6h11eVjVc=
//pragma protect end_digest_block
//pragma protect data_block
J/H73L7D8QD6g3Y+NYuO614/AL3MNiBEHl8azHbpaKfPLQ9PdRIcn4sJ1RqR6nrp
hmic7qDS8IGS4kO1FrIEIGmXKNJqaLyMqSyNUs0e/NEKangvJj5bkIBrdz9r+i6P
TBbHxVBAqxJIBEfQ0nq/LMp2iKHrzlWtldvU80bELlwi28OnAxoX1WWnxilItFji
Xc/T4n6PXDZY+KZo8iKKn3Rfk8r9ot5fSbPlfyasCmzzsF0MpjU6UVexcRTgFUCm
LlHsdK9Ti86VXo2mjzehBpq/uG8FGN2AOpn0RDe+plfRmcVcQuI84LIpwKQOAKjg
Dx0DzF6HyiM+IaPXht9TDw==
//pragma protect end_data_block
//pragma protect digest_block
vWhwohGD0cOASqVAGDVuYCmSZPs=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AvN8e9vLvVjr2FLnDxbtEgShnjHK79klbFsWKCyVOwQfjJU1OaFUwvvzfNfvbj24
tKYS9CzUppYEdce2rKy422Mo2OcutvIl8j/KyPOqm70QM4ACTtqQ6MIdgRjrsyQQ
dq1yS4IsRtIJQj0pJSXk4XjCGUrGlcvCGDiAc1nsAfZXHy98fIUppiJPNl3nvTGm
hCzsR/XjCvtQHWfUdo/oq2G6BvHoLANR5gekbqI70wjrLOOaZUc/HMzho9pwjLth
X+72o03ab5G+wjfOSegcKbv3F1I2BaY7XLI3PTejJhm/ra1dL5v9bFM2ud0lknm/
m6unshRD3Ivcc4msEFZ2Ug==
//pragma protect end_key_block
//pragma protect digest_block
V0Zn8mmA7dKadjO85F0X6pkZH3I=
//pragma protect end_digest_block
//pragma protect data_block
avsc1a0ZabUvLaAmB/SgGEw1BN/obXu32nNgwuGNG9QfcvFYRXTRD3cr4wQT9XiA
5+Of0JxTzaalzISlLwqyxNgzGLmOr+Hut78LHjJhKAjtsrkVrIDzSPBlYwHL1Uf/
tS69Jw/gf6mkgGH3+hap0+0qGV4EU+Rz3kBei1E3Ud6+y/EW71Y2RS4uT88rkAdO
sSE7mDZdD16/JN4KPzSGIW0SMQEI8oacATderf1mrxn3/Uk54rEn1uPRSUJ2efXz
zjGm4IdU3kdsyBqL8/K5A5w4A+9dvQQ6a3gf9gi0HRfyFMASD6MmRXy6aH9BqZxB
SCgrvSkFohgAihNsrnI3Ig==
//pragma protect end_data_block
//pragma protect digest_block
Iq2CVlor74XDmdVS7nqht8Mg5sk=
//pragma protect end_digest_block
//pragma protect end_protected
