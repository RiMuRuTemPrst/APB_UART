//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AZPYc547bvgZ9rP3TKI+ZPQ3j7r/T/eOLeuAUvYWlt5XJ1syJzYWMlcGGfb7/aiO
wZTKUA+6DfaEK3wdmgjAyWGT7WoedvOwl1kyFRDWynLbjLPPYNSR8mFvB67EWzuy
f8T8trl5ApCv1MjWB9NjEkcSnP10OF5KtvgG5/YfBSho7vBbrJkXFYeb0YUV1j9E
nnPGZDt8oMd+dZ1CCsBuC3sVWNmzJIRevyQRC60FTMRW5dfZiB9ZDa3w4uF3HuvN
8hLJJJGqidukQx7pGsBXOTXLNCVekklp/oRk6UbCIGmTyt3tGJLl3OwMGBgUN35b
iU3H+hXb6OBDCjxS9Optag==
//pragma protect end_key_block
//pragma protect digest_block
TN3DKA/rzBqSAtdhUricYw+OoDo=
//pragma protect end_digest_block
//pragma protect data_block
6PEAM6pAsewmdGdzFEfKEVqSWa38F9TLIBs3AZkR852cVCsODRRbVhBuscaDc4ul
epnvovGZUWCj84tVTIp4ymdy39h+ps8DDQAEuL8Ps4wdLRsIbUUiKThRvP5nPUt8
7JWyV+kPEJ3rmzxcM8V/n+zOQq8KXwbpKbehHoM0fPs6R133zmmezvep0nI3Cgz4
4YINc6+s8QI4bQ8CotB77ro6GJqm7jwX2nmxNi+0cwdO4GM854VoOYyYkCuEr0Eg
C6yDHIRc2uoHn4ncx/Px4LMDNgv6O8aHNXzoV8hUwmYRosb/F9AhFyekoh9ROXbs
lVwU78A1kT2Q3b0/FDiqZw==
//pragma protect end_data_block
//pragma protect digest_block
WQ6hBP0id1f9h+Yx1N2wE5AQdHQ=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AP5wlwyAZ+SQeM7GmlRhOJFgNSAduJl3V1UAu7w3ZvbC1n64d1hFp61bLo9cgy+q
j6ENECeN4/52gftjaccOPJm+gFGifEEJHuU9PDWGRqA1qOrnCtvJQKRSXdRvTChO
rusKdyCHdRcpv9TT26AsJRZgU553K4WSh9tCe/ZuDhlbXwVTZcjwTCW0U/MQjbV0
xseJD7QgEIp3eqTxQoEa4nzbuT22Dgxe71XG1W+GdKgGSzz/TBG8A3uRJJWbOUuq
BAbCfFKUqcTY+sW4lGm0KdN3IbkHeYGGWq665U60w6Ie+SISc1HI+pawUbr6qTqq
1/X7uSkGCxP+za7FgWeIsg==
//pragma protect end_key_block
//pragma protect digest_block
VbiD5/ShLMjCrwrTjNAdl9V3XnM=
//pragma protect end_digest_block
//pragma protect data_block
naBYOWahZ4IsL/UVItKievtrivrpbNjTC63mE6bVymamG9Zuy8DFrErVDSWAhzyh
2NNoF+JXeIOWbo+gDcHbmcwHrK+mB6ggztu1k3636Cb9rG6LwmxLM+1z/aolTk6q
HeTiH6kbwxPq3kQLw3D8cS21Bsh+Z92C8kltbKjVu1SL0/WOH3iCYV1y9SXEtK6y
RfOo5rBwO2Y/m4p+mud/0C8EtX9X/cK7bCAmIcy1TMsyHd8RrO4f+BKCN3DR0bzY
nYl7CaIni2cHkPr2EtJQyJw1paSSMmnpjcK2FsXDaasfsNWBmtTIX4Pxan8vzrtu
cQd1GDM1YsEUmTlKqFp1pw==
//pragma protect end_data_block
//pragma protect digest_block
JVcE7piHbbHgzXNB4dYefVbBqrM=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
ABoyxw3O0c3KhPSDADz6ridcExRLEXVzdp7b1ORyJfPiMK9uYtA7US6sYbjg9csi
Ktt/2xFz1WQ1beZv7Zgc2A/0tNbZRtqZjbVP7RktXGbZiYgdyGec01orHBnqMhma
A5jZAsPHh83PvB0MNuI84Y8bTHnb/ZznEd0wrilrVb/swki1s1CSbAfo6Eovccz+
6zYdAZLIpQU/1t7rofNgLuhORH1ngc4bKOr20SmT16xbj4vMsCfmcdF2pM5ukac4
VgXDp1DuqBG0HpqNYTejp10sYaH53dmTtaOq+aC88klfSlRuN77u4DC3HiNLYNMj
HbaOOhUasFFgc2dtd9jzxw==
//pragma protect end_key_block
//pragma protect digest_block
BjiDJnCF2qmsWxufqPpiXPbNOXY=
//pragma protect end_digest_block
//pragma protect data_block
kUPbPrFZItI1KVWQ1USTt5jqpxEMDgc6qf1utQUsfnzRr3h6+IM9FDxygSTJr/WU
M6wONkjHf1MfXQf1iN8nAr9FP8TJbI7YeT/0UC1ePBGaVhUwYt7Kb6bbynF4t5Os
YJVGw6Yu6hzw/E/LZw4JJdIsoM7OGYOTerDwpXSzdPEuPMzGZyNcT2RWcMqVefGA
au13rY6GnQ4pwiMPlukNrwM3v4u7frWJuLkOSaZ1S3c2dQ8qoNo1FyOdHFwqtT4q
EN3jj6Js/xWkVPL68HqJFTBzm1cCRf/uGFkGGeY85ieNe9oIcYuK3Dp2OVeWtSa2
nY0RmI+T19igW9UZZWdtcw==
//pragma protect end_data_block
//pragma protect digest_block
Wf4sETJlAQfiiyBOMWuZoY0g5xw=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AunKWw6FxfXZImQKg0pg9mdTJiLBsYEDW3TNbrRHro4nlUwtMJ3BtCBp/u/lp4hm
Oyjpe21RKA46rMUuxYlim1HEl8vajoE9vyIBnGLjsw1JWUF0ju0NvDanhr9ug5a3
xJCSkNrZyKbkw/VRfpn+Os8+xUWgjNVpzdo0qR95/atMVnQaI79cD797/P29TSyB
Mpg5z9CFLz2FvP3CJ7p7TZiGEuFgHWUATr6rlTkRGx0TiIjJmYKCAby9m1ILacPn
ptf1Wl3oEYkPoUKh97ZIMaeFv7IwmQ+Yr8zSxsmN4dXBZEZLGMtv+rr8Y3zTWXhm
EE+9NHncnUYTKS7SyKTZQA==
//pragma protect end_key_block
//pragma protect digest_block
N8td8ZIGs/q5qFXZE9NPf9An01s=
//pragma protect end_digest_block
//pragma protect data_block
MmET6S6VVIRSTUBImeUOrNMD4XVZW4Jy7ctf+KdNPEF6Ec2oujniKXnhUL4Vxy3u
X+OBsek4YPFnSkCRjXbNEhCuA+w+Dr2hnagXmQ9uTiCjdaJXnulKfYikO76Q23wZ
/tLRCxmcyer3AhQnvhlwwsKAlXx+7hweIdrRtiFR04unOr1Xo/FPucj4Uq/qLBvL
tTMusKd5zDFlPUhGuOfjZTnNnjiDt6LBwdWHwchMsz2VMpaZxxacwW5VqZ3NIUUD
7a9VJqZYs/P+doox3arqVWeJJ0UX4ql4VrxT1c+GAuCopR/sOIC87j+He54TVIFo
TgBdDExBAkfQrajipY8iSP3m01UHGIDPFhCoGiFT0bZ+zKtKzPVH81Frf+ZoM31Y
mav61r01hm2H+VieJJZgvpK6LC54EVUluJpQSkKflimFrRdk7z8mstx0+OnKLvb0
7XUIvH79HqVjxZN7vxwNFsYU/Gz/sFWZJjMI76cc8wdMmpyOHyt74EG1yxi+jX6k
EQJchb71oQD0aiFSechktYTrgC3s1220xCsuh4vjbiNg3ZoZye8m98UGQ/OAWRkj
HFpk9zqkBcdMWr+K01UuQyGsTVd4vKiJ7jRG9LzihKeSzE6l4OecG4wYX9AqfcAj
La6ZQhF6CFRo8ny/UhlF54JrfMoCuJb6agZOdBj8VWzokZmOMBjetI10Gm/96586
eH2PIchYx83TBoDb2gdK6Y1SM9fdUxMVkzPn0Et7ZaqQCEsNo5J0VE4HsBPIObVN
vdW8bmIhE5gbRfcRYQ3gZtybUIXGD5YzLeBQu11gY88TXmu3yMDGgtNdoNOhK4Pj
hpi+pUIxn9yZoygj5aA8VBCy6pNuI5murOufdenh8hKSd3VK5U9muOi6CNmTE4xi
88H2T+/kSxCP6dlcXDVYeD8gSVswPCihVnHgXfo19b3fSlU/nekl9uPWM224lH5e
2pi+HnNurUIiJMMrNKvRYc1SltnKbk7oDVs7ShXgKd7AV07jqi2p3phqWhS9hM2S
nadpxCiEMTAsPWntUv2AVV8wyi/VmNVzah6anDrqGc4vqVvw0DVuSAAQehDFOxL0
yL2bi6exhhhToVYup1iULGpLvsyglDAnK6Nc/MFsVv49tAk+q3HkozivKd6bDv3w
d+asUCthI0BrMS6KaSQTXBwpUdZ+lWiQDD6MvgI7lXH/kBuCC/b2oxZFstYHOLBV
pCvCtWlXYmHtBhx2AxUNsw/y7knhQCHRnEvYkSs9k3Jrz+YhhKWrmEqFjoEi7QDp
hMTZ79eRiRsk4XNmrm3Jr556TaATwuYeMnrfddLJv31EtIom3posUKTmD7XcAe8U
D0LTK2OAtpwcrig36KuBtyCcs4S/6P13W5FbDzzKb5K+xtlYEVMlMP+5F3digwUJ
iro0rVMYrMJuwz3pMgDKBMj2EX51vJd/1i+QZngO4TIQpPlrKH4yx+cacKbJG3es
IQvIwYRDACMajoKblBzDLuczAcTjkpYziuriPa5ormidHi4ajTmkI4jaXKqGhdPv
hmmAKVI0cxlWODf5xqJOn4fYXdybwMut0oqEqa2NB16tELVApUru/IUXL2Xcr5Gq
F0rssWQh092Hl+7Y14XpKICUss+k0a3WI5uO+GLuSLyrfYMje5iZOkEmUQpGot/P
ZzMJXk+ndoXTBel7Z8tmy+hEUbqaQ4S9JYgRgRqfCfoG2ZvB0GdNhvfZqEaadfK7
HTh4fJXSI+oJJM5NmVVToHynBEtsuS5fxMBY9TMz9RzH/e/Al3CqZjCttk4oQfyJ
F2rKYcxVDliK4JCh5nucGSjRUd+XeboK5qN1po9H149A8FHA4mQyvXe+OR5mu9Zb
NMb2zQpd0XaAn4Bp09uewR3eanoqfW7z41o3rCQ324ic2RjvIi3RVCjeAmTV9sIU
d9183dkVMlZBanODvEyjhHkG0f9Z2MMComVjwbNcczeBTs983L81TrJPk5uTBV/Z
jMbeXIx3KJ9xpTUqH4v9XIhlWtkd6iba2xuYP12fO4yBD0E3vPs4drDbiJCvckhs
TAYktcvLWqwUmS+KdRA5iXydAaNR5avoVW8lzd/Qs//PRlthRzQ71abOGL5GjIyo
NORXZy811x1Y2qn2ionggKVZWmTETAwcRTu51t6qkk7q99LgM8yd1A0A3H2fyaD9
CxbX3Ho4GYgz7HpIRRCBDg4ryKelSE7w+bxMp/+dQ1hUyhuxUkwX95OyIRhhagn1
mXEFh2TxQ3jvc3YHxUYazhMaz/NLSdppSC4Yw8KuUEK7VdG/aMkenWlm/yCsRtS8
lyKcOb4B1Y7h7+Z3mvzkwRamvNiAegJCmlEHwz7YctcCS3FuvBGc9ZQ0VtkMsTDE
Omf+0xLHXs/mOJhHN9zuohyHuKT80bd7qltyjBV/KnApIGNR0bP97taRIwtz5cy7
Bw0FsyiW04D378exRouiuyuQl466yD+77V2fyugDzF/P+dl30yrd4jTs255fW4T8
cDGTvS3+PDd79A6CzgRhdkTAA9qmIT9nAM/JVpg7eN1eKdSWM8nd6Qv0O9W0eGxD
Dk3ixOlAgggiomhNFUbYCfRJU1TnFwNKp9F+5MpTe1j5LjfTf9JUXZRYKg99WNu6
ornd9y2pCO7fhS/0SppMhigROv6XQ0urZwSn2ptSysxap2TF53gW+UCo5xEbbyE2
49q3iYkIu+3bekc4ykHKE8pi31rPMS4Nua5vBk3ThoZxBX6q+3aHqt3FRmacZOUk
j8c5LdH0KM968t5PwgWcFB5UiHfOGTd23zkssILxUdfrDhfviO5ERvDfsaKILWYT
LymS2i7XLcemsOep6euMgdoaRjDMcj6S8JouSapmrR7y1wasx1JyT1hzDesW+oj4
6JKOAvhgtpcUIRpR/9KH4n9APBRw18yBtgiJabDGtnCMS5io5jfy16q+Jm1fykoq
6117btBQgvmdaVeCrCuu94uhOeLmaOBy/aIQ2gySJsLhLIB+0YTjJf5KVmz6Zoob
gBTTeWejfDUgaO7i8PF3AitU1/ZInD5o89+K9b7fy6ou0H5n/QBcVthcFHsNVaf0
/INCDhaqPPIK0tvRAKCEFPk6heUlz6ChOu5sv+frcA1LCg5XRNHW/zj9PiODXzJj
b9fhBXGRV377hoT0iZdtbz5AEgH6ic4yheG9CVe3rSS2nQkgxKcraAoCCMoKTDp3
ryQWfZilwVwoTHG7ttFRFO4pXL+tJwYZYvRe5zbfbXDYUDoU3z/HVDXksm6PSUFn
ZSImJgTXuGJW0FbveAfhLsnT88N+q2CFRF9IrOVWwc6nGN2ytsJteXJhYqGv9NPZ
fns3h2ic5QaRl/0yRZvnH5jFksMqll3bMcXHGAcqIqUcE241g3GytU4GTOwg58nO
rCaFsX7e75wvqhehiV/Nhm51IYAQW+N4zoxSXoYphgGUA9N6MTKhiZO7Ut9IuPJ+
K2LcJRFyP4U0UcCf8H7UOaUmuA9l3H80KM8680XOBSBDP37GbX/YfeD3sq7Q5Q+4
hqSVCa/kaTLKA6eKgWcIGEAM3k3BysXqVTghXRARYyNjQ+8/8HnatlfyDaALDIsM
k0owoP8acLtIyWe6t6gIm+vlYYZnKK7FHoTyZUleC7/h3jJ98V2vEq/rTzHpMxGj
WZAx2oyfUz9VqE+xq1rIURSIcagfktnC4B8/DJoQ9WYpuFyeJb9CwT1zLQKxn4b7
YbMzFlBXNvvipJn9m0sOjMoRHMBiwKK0jhYc07tfKpSNhLzE5ECxHtCr/CqUMd8x
KbI1dypYRrVoMR1gKOP5Ee6nvGcKPG/+GYYI8cqRqy0x6sBiRo/7fRFvBzPHea74
+WL6qyVStP+7+NpfkdDZgv3jDVoNKbZ/Zyaz8W92oyKw61F8ZSYHnoHyl3KJF7FV
B6GtE+vBeTuEt7Y2czUS5aVdOPYhMtxv7hKAEXbZ6gfDCbpGtfYWnQXnLcS4XgYq
jHoTPWRlMiPWYOM++fQJwi+N73z8tN6WHBY7D6OcqETxH1DbCrEf9ag+xD37idsa
yl4UIsDF2AhZaOlYofZGczUVEPa4k3J/3CAcOCPhub2iXZyb1+RzQ4wwoZm4Rt5E
98LOd+FMgM45fKYPXziwXQeZTkHgbPps19ygZruqY5t2t8xoyY/sSj10a1/hSlxs
v/yck0ugLEvRJegMvljOMLY5euZ6cITSWcNfTX9+HjbCLO52ldoloIl74r8DApPZ
zWfBjJg0mafhpLdv0N8ofJu1yVliLRFuIpVJqMY/W+aG4t6FehBtP/Lmtw4/MwLz
LKSNbH530jK07wJImWT4DnrUarIJsnJNO1KuhYdTRY/Hfks+rNzWYLLM4CVD0gvB
CfQpXWurTMM1Rv0T6+KFXDdIBZu4LeUJnEX+bDdzEbgJ0/9D0i6nVUfVgCkk55Go
LV9vZTiQkvLPlsOB92B18S0xQnBIiU4kFE146Jqy3RMIfI+a94waJvXJKIwTbkUb
6pTM/BE6XOnqPfago5jVgLESCdflYrVchw7U1PIAMpQikp0c/pkIR91k8e/epaTn
FMkCcNjjxUZ57bJyauITSMUDMPNFKmKdzvHtMlmpPDvkj2O66HWcvmwbcz6EKg7Q
2R9CoyxQjRutqndN/dUWEPmvawDXl93GZTSH79G3LizyrSLKY1hiihGebwsdHP/6
T24Wiv+lje/PDjA9rG2446jnV61Im9CMJbrfFvctY1yyReiTHsw1ps1wUkUEOVUQ
63l9e5jNACXPOQvieGcVoL2A/vZBn9RJXU0hiHctli1x1MQq/9ZLdTuVe2EHDDd9
U+EVx7mGDgcd+DbIi0hTU47jtNH4rujxobw1hgSPh8RmN/5Y81dyRC/IdBX/1bG6
slw11ixyIWJTJOWM3e/SeTG7SVDcnwCSUNN6/p8/hkeG8a/LS3thqZZTUCd9+z1j
bUJDacUXVFfzL9/tKQG/+XvJok+mAh1VjnNBX8Q7t2giHMEDYe2DggMZytA1tIw3
Tc2qypuSat2/raxF4LkA34r0OLn8/pxyyZEw81vjg78v0qjkbBJRcTXpZc+66z7M
4POBenqTRfYFFIoj0wXpgJr8IJ586j3FfeI9hy6E0Tb+ph89L5b8Vvh89fr/tJKy
UeIB1RCJcpf/IPYUicKv1Yht0hgbAERU1Q4W4rh7YUzmNNPiBLmGUTB8K4dLkA/3
tRaIj/BMBNmLEw71Cu/mNQqNekn+UbyYxeV7pgmjhtGxyyxgbm4yejUMmLmZQKvP
EhaCeFCiYicSxmhaCDwuk+u8DNK+I/G4MBZhmHS1jJ8kf9HJJz+oqrthI19yCWP6
W+uwBefqr5vuzCyQqSQxCo9JL/7BhFfg/tdgfjyhJNx/PhpcWPSH6lbBEspRmWFu
aXXGWVQjWxEg9GIrkIeZ322tdoIvZGqA4rRFtJeDfyswBZUoqDk729ze0OUnBAj5
QG7tuutNuDYFY71YngOpJN0pZ456jXuveFu0K/t0D2xsd7hNP3DS4nK+Aa1ran7/
f63UM9Wxp8e/Q3eARU55Z6WDSnahsnP/oGulQEjyVnJRkguaNFDG1weapEcYwIMI
cOh1+M/adiKPmY7hsN2t3w2dqeOxkimABLDcEE8SrxntRGzYqk1wi/hHBWWFnA5A
5khfIhZcLjOp+q8TDeVvgAfUSw32g+UZePG0xMCXaUQn95dpVWI+NIAm28lL0U0m
bSFC4Oak6dQDOQjSYQkr6kdByzm2hYg3WYLD2d8rZlFjmVtwZZr5x3T56WE3dTiU
1DH7r79X4MY94TT+mJNGjQ4XoKgKon3Y4XYDP1xYK3ewfd+e+D4KX8qIknx6f6Jf
LirYRcklyE8D+YcLf8HSSz77SlvCo4F74HxDcVMrLNZ3ZqWvbsIfgGFcWqrQP0aG
I7c+yDsbO0M0KgOk/gWln49pmBefBc4TRN5lcwg7LwH2Y/lRi9MZoHu+RLkPyX8v
eMo5cUykw37s5t/a4qy/OxTn+LZov1YdH358ftk3E7jl2y/k/qudhWyCyM5DVjPG
PbjxwzNAhwwI4VBViigxqjhTuEMso1v2eXi7+n5V2Q2Rux49Z3f9L8ckAH+//RZb
VYc+8KGpmsZFvTsinXVM/WNhUbo1ppwCPBJHM+3yXIGXR5v5LWiXmyHMTsL3mKP7
PnQW85elUUrWG/YGEJIlVBleFCekl0qSqfyr9ZpsuZwJfGknOEdrmgWvjKw7oyz2
8Z60HNkZ9+XQbVl544cJsYx6uxUNflyyQRHQd7GQ5yWN2DLp8CMih3cDwA0WhFBe
j2766wCERIKHUIQESD2LyZjyHzktod8dDGlluFBjaEa2trdNGoiptMnOXaWYIgy5
TveQOXypPJf92FxbPYH+3AkCAsL/anLMi4H53z/DU/7nDd1rgguKn+AGO/3x934k
hGfb6C4yXcms6RSPOqyzUZ3klS3OwJJh/U45DIiDVn9wZ5gk9wvuMpf/KN2QrnMG
nWV2XU109BcNusjXZn/nvB7H1lpH4zjCWwrMOpZG9sylCeXc5YRAUWLghtFol9ha
/QSMZoagS3e06596WpkeKXZluFt1MrhPUq8qCcOhMFNEOtBGniq02jYRcc7KVZ4/
edzKmWVWigp7Rhaz/AB0BpX5KKuQflsmURrji4jYcK/P/nKiRILrht8QXivud4cJ
6eTFsjcwZA0+tCcwstOogMFR/WCSUFy28H+ylbpLq58UJtAYrulD04YagqZMr9si
MmIfS5ExWM5JxFtn+CTUj+jRcJE3nnsGtZj0D1WD9HCYF+weIkmeaBlTFsyn7WGU
8LFjSGV9FjnI93emzp5lS4n86/DXO8//PQdEsz8T2rz45R7Zn9hHZro30cqxfjLv
IDft++btCUZah6Ks3CwN3BBjC+Uod5HdEjmZ15xO9YydgPYoJSiOGQU7GTiU1nOK
C5mBk+OLZstt+jCyTa1ZNyMBrQeKnNZmCrlxeNSxAmAvlDHS4nFv8UMkW6acIHU5
fBwuJxbA52VgkbjRrozQ7wnWIFe4Lr065NE8J4yoIV4COuw7QaVq/4qSYXpxIi6X
wEbdf5wQrTKINcYt00YVQYtvOy7I/VQTLwFT2hSC4Z2B+e+cbEAGHHszSwWN3qYD
SPHga6OUfD5mVS+PrXVz0p0+ISSVA0INXLRzOU5bWKNHb0asm9YrPuBHfJwNAkF4
BWrNy+Uyp+O7xLVMEQ/pR40FCLLuIwo/M9hRMBkWPOZfGAJgVm8xir1BEk0T7VSy
W4V/rJWKp9UFNaBeTPH3ew7XLgIV+9jZIpIYxFs7q9s7DlEsCcpwp337kcs2qRQY
23ofuyw85OVpEyWAZex2uCIjfD6tqD70++Jr2qKPHEmx+B5CGnHnQMokJG2EytLh
izEUCpPsnW9pmV+Eu8PVEg9iihuvwOkp6A1PhBIkAckfGAoqm518i8YJV/iApWa9
4UoLBEfpk9+12KXzqTNdBktl37TEUwcdIYkT2ygvP5VhTPv9KGrXs0Wr/JQAATF/
poSOlcxuO5X0ZrIKDTQsuoJV43gjMZOwQAVGRRs5uug/gCcUfhC+wptbbxvGQkFQ
87EpFqMRlMV9J/KP151+uuX2QlJaTnT9M2mM6vf1x8mSyxq7RJNc1oNoSIHInQhp
BvOs/UWlqzrDO7n4HPS1+1GXqfRl6oVmXQYnodgCRjW7uQ/FOKoz6EpyyFtL1Kel
qzR2CZ5N1KKWbAw6PMjb7CAEQya1VV4f3IW/pWcTzwpQNs74dg7pLxkMmBjBWQ2I
cWVu5V20a+y7kqoQuK62IaeGu+Y/mBcLY5s3FZtrJXHgS5yloHpEDEoTMncBJwK0
nq5TyIJYA9S/cva5jdxwg6Z79DeyNx5bcTLUw5WXIlRh8NaxoQ29q7ppIl8hOydb
Htf2iKC/YjaXEkTIPAETCKjDr1+HuVNk9Ag55Tx1bNrHiibiFVqniOjz2jYgcNEt
99ZDYAFECqziUWF15OIxpR8dcCnOHJpHErMkVEbXNIl7jhcawCOaUBsIhbmp5bnC
q6aT1gQWcGG4F7lKE+S5Dl0T7x8vGuEJpW4uS0iu7H0r0flFUof4Nv1YNVrTpfvw
KXK2eNP1ALJY5a3MDTWNC7kbW23zcfA+1yFKgWhcl/IE1ZR9Trh1rz7UNfGIZTW/
0DvIduY7Wcjm89VCsGAfZjoJDn6g4UkVvySNGROcTsscj1dMBlUvfT7ZKtPn8GnP
H4IfcvJNgDAOf6BcEzZQ+kaEXVOkTYn6i1cEfeYmHiwzj42xK1eS6CTHGf+7XJet
ah3PJqjYsiMGHMLNJxNUsIkXHVFpdJvb+JyHGqwMTgsyd4UzZpO+Va+6LrDAMWWo
2nJISecjW5U7O40SXXHgDA2r0ORoRomjYC+WI7OROWBScB3vLVHGY600oOVaT6po
h52vN0kOuQm/OhkzN87iVct2wL/HWy4cAy1I4aDydB5iLJhqSplYwNw0xX/hbCvn
/BemfTla44S/fV64+Qj3HaZQ5AlLYxcdLdDwzvR+aSx3HPW+NvK7EDhIvWBFqFT8
sKpDHUgu1EpmMBH7IXThKOPKqpRO1OtfX0bzpJ9Sy/WkCkxVlslQb469m0l5959+
SajQpFvFmCU3+V3pk5mDn2gcvqjFTko5rsl2UtJ6MFV6JhzLkLsUYQdt1o8IpgW3
AAk313us9jfihC6TYQovsArx5qGotrxpJsnc4WBH7tUvfWcrO9xmSbfg8Ig0/O9a
gpqwAhhhe4GbYA9WtKNTsOGOIOTWRPX7vV45o1Vq/CG0feNFnoyThZ1bx/ntjPh4
XFcoKxTs8S5IAkAjtkTx3XBkFhYSDoJaMPGd4dk4xNBWkKuZuyE+W41Wcp9TlrSi
qjB9cELfMG5zCHoZRheDS6fU2j1MXSj5SuwGS+gVjuevgVOg3xLoMMPa8wL7wEYn
SGHxYZzkiJGzCBocTJ6fiI4UIUsk7MqIH4YDlzDGtP71zM4qiFx9b4OXFt0DerZB
G/AerFwYgTNkKmTB/wWQ9wM4/csuxD6OAmzWZ0a3qDiQEbnmC1VEoZfLtvj+5y36
u1uQi/+bVeqZEZzyuUaAwZ692kgFVBeE9j7m7epS8cL28qXtILXScRkzNE7ivtZ0
ZAS2dlXg7Afjh7FxLD1k35CIFnNEQdQAPSfuuKGC8cAslvgT9WjfEo6aiBGeJBiZ
KkDQRFY6VI2QosMeNzKmNj+Pj6o8/ObioQSCfKkh2r8KubQ6kxnqai+SrDWahmTQ
1cSNg/JlyApBwo63BwtBL1kv0qgCaS0pseAwTnwLdN2KtPsS8J3and9Ma9+xWXEF
dwhlF3Hq58ptx7RNTlUffctRZ8+VOwHejBfamACRME/yj0x/6WvtlFMGhSrLtEm7
iCxLnliha+KPuD+GKvQYaHa5qb2ccSYPisKUc8cxFSDLJ2N6nvchP1WRnIAbUnHw
rGTW5aQT3aD7bzIXmvkFNy6hrOiakhSgNf8HcN2tqf70xggezddVc5zHWIsA0mQb
x1ZTU26cHDdn+nUqRnBWIn/cI6k+cFmhHbibj+k836B7SZXqLmX45P2L/VMQWXAY
cE8wEOw6esKx15Ep7UALWoQFYkT1YxxJE9O66RLh1TBCrrKggUXjL77FG5E99i6A
GGcONz+j+Shd13VVMNnJ/zaGZNaiLP2D9N8dpVu60DGvxRuBi1F3btNMIJiikf/l
Wv4fqX9tXCVAXev/zePrDn2WY/PkdeHrcjx4PH0Bik7Ea7ADBNFIiZv34ji38mGv
NB4fWAxQVsMxFMYO8RefwKVV8y+zpcDkuFSGpQVlvjj2Pt83osD7WoB9z7SXkcrb
kCGNfTeYk/gShzvc/0PKlUU7th+xWG6a29zAhXL/uF7DNEcWbe3TWDcnLCz89zYC
/+s9poeOs3AmtRunbsrLKkbtaGxEgJCfqPI2Oov2tLgjkfkrfroslqSiu0oDvNUD
0AKf6jUMCwGDZYrF8jbcqpRcGxdXOC4C0suMW3IIU6QPau1ZLDj99pydEy+dVtzQ
N3TUvtio9CMy5VIZXL6Jls+eDnx05Yt23xVqoeEJCq51aFTP3UuK7HWhwLiL8Rh3
nkDZptQC7YPQ/AlBmk3lfd65pLrkHuCXjVqnWSfX/hgBpZUPRHlXDXERQKBpIRiQ
HlE9WI1zAtyBX1L462uzTxE5M7x4RSHhAwwCtrdmy35K3BdD72GZrXczBJd1VH6X
HJRGqg3OZZDpOok9itE7DyCxfg8xXlBqkvWncWc+cYrXGIdhzB5PncYiP90d+us2
KhvcHjxq7ZTYG5YVD5SRmOt99HdtMUl32ytJZlmiqvL3aM8dmghJ9dV6BZUI1wOi
I4sVRbavR7+TvbdP54ki4v8XZe0H/gejfE9tA1ZmSzkMtijJXKHbUkmtxlQS8eqp
hL/MeP8HZicW0+Sc/fnORoMWMPMsi1cNRS7K6Upv5/0voZdcQaws0bBbEXAH8ekb
CB7QuO6LN6qYVE3v0/UIl9z1mOZkAMZVpjESUwVQ97o5bqJ7iq8w2o10PBk7eZiI
kDxwyNtbiLce4I+xXYsrow6hm7MvcEiEFhQrxZuEGitkcSxi/cGI5lHfI9XKuDdB
rzN53mquEsBBwdtQ2kCLB4nySW+5eAtInTdkpHgeYnj0yq1siz38A6jr+QsPlJ9+
MiNYBN+Yb2xCar02GA74i6kHijbq5b09ZnqRgiFzN8QlHToY1ZPgwozjmkzQgrxH
y5lY+NokTfe/Zga2yIVQxaJEgheOUbdh9nJg2IFUkJSAiJn5NsMfsQgvCB1+anjz
hwjoBj1MTVLmnPhKJM3r1WpRuACFS1oNaEQw78wYfHed5NbQfofIjQlTb5Ool7os
uDjyXH9n6srFovubz4uS/dueo0wW++2e7cxsUfB62kboBMM78oePLzV6pxnspLA5
cQi7Ow/Cckw4GmSrt7N87mW9A2g8jYv2wj8aILpBnEF4pnsAKiOe9IGNLYN04Ynn
LiHdhz+fvpgGa2oiRyfytVSbcbWU47/zcRhTCG+BAgzPHnE9/HA2Mr1YdZSWAFpI
g6BKAQD7FwqJz9fUoLjdWgWBsHEQJYpyrl5dvoQ/pq1yyR9ePsuXJ3L7pb/LKG1X
57ZBxkev02sKUYSxeethMy5nrQ1+RU6hiTw1UxWQVjs7D02QVi7brfF0qOt/CYuA
Vw9ha/vUA0+7MKDX7Y6tAH0bTU166vVFSROrdkWC4xgRlmjd7pQV/2z6t6kbk6IB
TJMHMrLY1CgLlnuwP7OzRdkyzvAl4isrEOw+6w4zi+OJYohdByKa918y325ycqqm
MMhqH1ZBtQGSNdSziFv6xs2elL6oSUkZgX+tmURilT0=
//pragma protect end_data_block
//pragma protect digest_block
K1TdFZClJnC7dzP1jWNJW9ghMCk=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
Aoz0p1/W7G+0BCbakQy1vDwBGcUz+aMz/HePTVSVSAVfLFMjs7XXaSMn0ipoQEZT
CeAjbjy0QLSPfNZGYlBqmxYn4xfq/dNQ2Fae0vdJFHQxJw3s2lA7e+JNcfEpnONP
mbf8Ne4GlMMWY0XKU6gtjbBoTdHTq+44lZdLrGATyRCneldPM69UR1CXQM9SB+pz
sLa/1ktMR4aly6/4ADNva/ko8brkw0gXVfhP5F/eu1jiAnkBGSwZG/zXaX7U/dP8
aQwdM3uZWVhDWrzR/BJqYn4Pl610JGErnJ+iCR1PKo0TtBh5vtOIRupfkUfbXPSv
kAbOBFGTT19xFKm/OfuMQg==
//pragma protect end_key_block
//pragma protect digest_block
nhIaIaQeySuw20khgQ72xb/uySU=
//pragma protect end_digest_block
//pragma protect data_block
FHnQt5ARr0NjlkW2qWVySkjK18FbwD5ZnxZCslPxjAAuBuV4IXDSyxOfJqg8TALe
iTuNnrRckiFSW6M1XaNs+F92jVrYxIyyLJS7bditwTqdt4oBTyY5nD1dFF5g3t+w
ciSRGnTD5AoesbOcL0bBaSaDJcALlfLaZfH4Y45+erN3pm097VbovSgNKifOfQRZ
Z6yTdAMyPZCyaO3My4pkklV30gGwpZso7JcEhgKFIvQGaWNw1pPxQmQ0zRwT3u4J
N5POqlSCqcpDfx0ON3NjD3+PwOkZ/GOgm2449hAQo2N4ejv2VGzyFwSSxxNdxFP6
kFXLA/xZUpoDwzoAjJE2lA==
//pragma protect end_data_block
//pragma protect digest_block
mFRlBbIBjmfBlc0v9EcAAXM/hGg=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AD+xcLkvXrs0gowlEJjjDKPw3ptjtcmqdWwcq9TzwqyQ8sUVTQ/TgID9Ev1bcrLh
hvj2fHzDiLZMMNpUOhouBUv0gmMBCO9xHpKFos7aglVEH9KYTvD88g9/TckkJgni
uXAp07pDeRQn+zVUe9YWM1Qv/w36+XyEO8ZrTSlHlQOlba+UW6L1gFR4DrD9ywE+
Yxxg9pzVA9evGpY553dV0QQk24boVFSiVEXiD26lhsIc3yOotD3j1uJeG+7pHvah
0ZnzOcBVlHUICGfYyqMLEjtoV5G5UcW3R86zZGuH6dKeWNIwl5YZ6VCDW+hjLQ71
hy8Z9Vuy59siEAkDpBdASg==
//pragma protect end_key_block
//pragma protect digest_block
dFdogoy4IluoscvUqYZm5MVRhrs=
//pragma protect end_digest_block
//pragma protect data_block
MoGFYui1astEzrpsL2riC/mz8c4Hf/4B6xnCM61EnaLkrObGM7mpvbwQ9mzLV3SG
7TcapkdEqgcp42bouonyPBQ7V61taGnt6mQJuMverXXfqg5kZLRbXNmUHsiaupMn
9SKlpkOxpXXg7tjJUogTgrg3hF33tHaoMp2Q/vEXlEXjznuU1j1Vu2CdgQdN2x+A
Ag3zD2A9gTymGhVLhWVw0PP8L9JH+X8m8+xw3lL610BIYoIDrIrtLN/lrDGGDjFq
lSUs2xpD1WD/PThDw3tPUhOfAmpKFf9FMOd/PA3qxRAfE5IDzrH19Fm5aLSoaodn
VN3ZVeD+xXdtO3xis30ZeQ==
//pragma protect end_data_block
//pragma protect digest_block
GYzfROHjNz2USiXDYDeS/u4IadY=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
ASUj3K0pbchSh2TjWzCcv6DukOk0ZmewWA1ZlkPxBwd6CfXoAiVdoWKh2KFX2wFy
QiDGGVENwbiyrsCteCxasBm85JgvaQNUuCDT0UhxHQNeO3hTfQY5ZtscB88cbMSu
Jf+/iI3MP5bNjsf5esVcOFa3nCzplVBy8VuXIKbpvYYf7S6DiF8QlHeAzV19MEZ6
cDlcnrVuQqDWd4iv+KpPLDSVlfn+YkMI7s2/Dp/xX1QG0VqStFdQxcrYrXjSf+Nd
4jwUG00jtXkGcWJZkPArPLSe3VsR8bh4oVJDZMnllKMbt6tJbtlsudnLq8myYXnE
61YUK/J8oEa+Yzy/ysVueQ==
//pragma protect end_key_block
//pragma protect digest_block
R/Dh2OZBwAHIRln6NtlQ7HBbQXQ=
//pragma protect end_digest_block
//pragma protect data_block
8aMr+Gzdz2LkqnYDZsL/VzZSWz2B27EOuBUEnbKZhSI3yk7VmHJoWbqFGrqq4hzd
SiyLrwW7KuYm/qOb1VFjyEkwO8qtm+1Ntitp/GYIrX6TFD7auCZsv35OLBxRPd8T
fxiPcb9afGu2EarUTDjnZEVSunMjCFD4b9HdsTBuDtHaO2P8iOI2Qp/Iim93ceiZ
t93hx2515QKGH7h1FOaasfGBlYhQslSKEGmpQCjgc+EXX0IrNikwpwe674EOBdcA
XWkFLl2EGK0sQ23+2dWergks5vte64C1+FYMFAS8EhqyUtyLZSPfT9jUgxAwZOMb
1h4gdgd2gr/coGZ0+/4m4A==
//pragma protect end_data_block
//pragma protect digest_block
jdFaN2U0jpWWAnrZtZE/BfX/Dro=
//pragma protect end_digest_block
//pragma protect end_protected
