//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
mxdOuuVpGY3McCdGmhLJmoZpqTegCsyTcQ4O2AyQicKcgZMVg2yVZeQXm4CVr/5D
W+NwVMD8RycWn7/3vEYV/5//nf23leEARCoOCtORoPoCF1EwP2/n2Kh/A+2MShSw
vkwj0QEuLujZDh7NS9d2cPw6iTjgZZtquh4kyED85ocQY4BvuTsidQ==
//pragma protect end_key_block
//pragma protect digest_block
jym9kb/dOp+Ldy7VnC3AJ/l8c9M=
//pragma protect end_digest_block
//pragma protect data_block
+31IgzqKs2M76umk4KZ4BT/Bc0udTPzmykNfYPaqejo7t7xC6fL0SV7KjSkhrl0s
nPWzL4CPOz/n7AYACRw6dRxh1kuQrsZU1WGRmXGidzVElKnuhngqnY/oq/YcxB5O
3ABqAY9xaaQFqvfhdG3NyyLgatms4LcBDZepxD0h6TLtmxCQ18HKfaXjEm78neP+
f+pBXyPY1LAjeeUpr2/W5BSZ9nyQPiOjq4ygGPzz82r9Wamwpo5s0UDj8I7KHKF+
Pea8yqSu8KJol6fa+WsA+OFVWfiiqtgFx0F/6aTzXduJQprzX4BzmJScHqcmURPX
wu0TSOMAhuRgq8EgS2GQgMD0HoguDmBQBI5/BHrTXktvPsUZaxN3Zq3+tSnRyWYy
UeIGHwPZy9ZHor2Li9i4nH5s0TRY8R4GagkdjbTkSmYKkg7U2x4qGoJZR/jvt4VO
jghlJyvkJ+rDryY8V7KNUQg2wGvOgl0Ku7IVS0Y6XsbCnUzpYoXEeC+pmPBVNMsR
ZSbg88JHf+VHBiYFNaxmlWP3PLAweN76yQnK5MNBgixIdN6INBksSa7cLfJxl/m/
iCoOrN9AgeMqu8sddHbGPwTCp58EsoIw2tIONFy9lChscC8mqL10QoTUYMTUr1IB
zeTTZtshPlIsbN/C8c3ymyVsZt1sdmru/YoEsBQnnN6CFNcd7Lvs+kRG62Djk3ui
Vl+JH6aUwQJs7om+eIMGav31m8HZc4nCI8kEnjwABgYCnjPd6lEsnZ4GVqQq14BV
QfarN3G8HY37IfRybLve15Ioj9AHsWLxCCBrKGd1KhmlsuUTHbXuJgkOqGASlY2H
5kmklQD1CNv1wcvxGYmfNn3zZpt68JN+xq/rXw/dTZ4sDD+/ExZ3V8g8HTn+QrlO
z3gxDGqX+akZ2MoVWgCPU11OKHRpDhESqwuRPQOtaETDq5b8dbVljDNQSIVheou8
HEilJdKr/kS7JkNsyKPeh59hVWYsIYsJ8GP64RdkErfW3As/h28JWgCR0b457RMg
LjEOd416LNYfDT2N7IiN/1jd2wn285CRgLohX8GogwSN4f+FDwNcAj/ztmVyooAk
BN9qCgkhQo3nCy4Tkj7k4wSnEdadWeOI0DB9I8F7SYObmCFDJ/XA7PFXcOtO+hP+
atRnltZrgYhzXqyYThw7HJE/DTEbcA44zMrkGS3A0AFOoCr7jzYVhp+643nrxhZ3
sjsUce4wfaMJp/hMuecC940DJ8QQGQX9qFsTu/Id2lp05mG5I/9rQponyiEOs5hB
GEo6WRsTriQ3T5vOx/NOY62vES861nnPQUmQQfbAcitjg0+0b/Zf5jnfMiJpq44j
8ImYl6crfL7+2OEDpYJe3if1+C7d0afjCYzUD2JJxpteyf8mFIVFnM5NdW3e79po
tjHlD70t/2rqmgcvwNlx6VQ5Y9AtfLnusVvVr6h0ObQJqGjRsCS5C7oSlWRD6gs2
DwDxBVM7nYa0wYvv5rKSxmWN69B419gOP9fKeAqnkFF1I3KDHKDlJxIa2tc2+HES
yPJVKybtV50L82n1jLym3GNC7KIN3UvoU29QN6PrqjorTZl4xs5Sa8yJynsH2dgZ
bgu/vmvanSlcNNW41rDE9kJdVXc+t9m3igi33u+AMZss2kdtYhbNSwCZKXEKnTN1
vkDWkD4Get/gKR6RWv/it5S24803ypeV7P00Qb1Z+O0shd7f7xvyVYHjas1fsRsw
N/Un5Vit9gKWvpIDrKQijLYzby95xvddIonVYB13cmaaSPyK1j5T2/Rh1LTwK/+m
dr1In0IK0JzWASB/6+R/BoCjue+PteKGiVfETMHlHvtxnLzx3pUdZR5+maA4iu6x
xog81WBmreNboFFfxz+wkRbC0CyDTJR2koRFlTIBT13ffEPHRRv0oNyz02k1aTSI
ibgPZN323hkQR0I5Vd80fUSBUrGnzyaoUaADiHh40iDVaWA4OS2Bk+ZCbUEFTwob
K22bBv49eX7LT59rr1D0w1pz/36IXDGOoJQYym5dxeVjbs/OXKjWOSJqQjwv68dc
tmHjGITSOUsJw54sdbC2I5L9KTcdYkQWwl+4oFR5T86r/6qXZhTPQ1P/v4fqBf1u
yChSPBQQ5x9juugmyqOKu/q4BHuyQ9CvRLNQEezP3dSp4qF+oPi3jQ5nbI6LdppR
V32sJ7rkpHeJjxiMGsEhbt8s9gXkiJpCql+1LK6qyjEgA1as8qOdv4ST9HNE37cc
F/33r9M15P2mDtYbaHD6ThDsnjAhmtiaIQiTY9LK5SuGVdV8PfFFbUn+N1/XYkxq
YlkAdpP9AQrpRCXR0ZBRSq7X0BCsXKLpV027Kb+Oqj2vDfOaiqDh2kuKykdyhIey
jcGlgXwrtkdBRmprrvp4x7LwtDGB0YLsPYL5ALqN164DTBTBk/fJjkqbrDlW/QUN
0oiFBJvfDC+UjKTka854en7p9yRvcavGjO29ykhI5c7+6k+B1jTBdQcCGz8qf4Vy
+j98XB6rtd/h/S+5bu2czBG0EbE/3HF7TXd6ZG9m/dlavpatTBqX5teusoqnpvk5
MJhDRlBIUeYp6GbE8Cr51+5QelUCbNZrQRx2kXXbLy5MpfP4MFSp6t70M0VcCN6v
lYVJjyAUFiaLdGT4VkuLXjY/oyORdngMgh80pHk92uGJF5UGudkVqZ8zVPEC+17d
jOHmPaiyF4eOxdv4Hl3MjDwXTrjRgKy7FLbIkMpK/EgbBNbK9bEACPW0gKR8O3JX
VOeUGMWI1z7dSFssoHdujZ0ZwfPoc4sKwUC2A8vR1cKuRWQ5HZ/bsfnP6iot+f5g
Az27fd5ou1B6Kttg6lXAq8rn9rRJ664secLgyddNmW1J9lawmcjiQmrqIjRGaQ3F
A73z+GPLiInCmbR87WsUdbX+lu4hKBUcfm00xbkAIxr/JGXFQiZywzevDiNfpt46
Yb6143HkYmdLKxC7P4ba9MR3291t8kggwsWPsQGcZ5P4JJsTwu3p5PH3qKcwtekp
rx+j331Ep/+yM05ek6sCLnhonAZXPJUUhGYCc63qqsAE4+fOl0Seo2ty85mZVFU8
+T3kevKHgp+OhNd2WXfd1v5gd1qjfoJrbxm8L+3cAXfkGOyu/r6ZdOderPw4aaBM
rFgiKmInCuj1NLtoRygCh9iJf5cq6fOdsELv4x8UYvODyINQdGJ3B2r4vOs2PpsZ
xKfj500lfVfWnyPCoLjg1lOP9HonGpRM4JjYql38Yo1uqjNOdIplNT93irTC5HLE
lkgX5VBU6sZ3NM0imgl5SS3xs+nAZdFdHTCHOCaxLTbdBzguJeNzjzzfO0iOowU2
M6npjUZ0CtFGqclZeZ+b+ac7/GN+64f4hhmDOXmkGNxm+ThhQ6NTQ0/0HwmCv/45
YiVTvzkX9l3nvd7cuZHTh18fTdIk3DrzswaW+gq0kJ0HJjzkGqfbgqoxt2oJbs0l
NNxOcZmCSLqB+0vv3mHir7wiNZOR3HAQe2cjTi/KgtvV8ucuAdrAxL99npkmLinX
ch1+ISHGJw1+3uUOHl7ZTWd0aa4Rg1LH4L6USXv3h77h0IFTGFRYqG5Jgw1dwb9q
ABMZ2MtGrK/h5pOFzcDsmyksc23f6EgcTYz8HHmE3CsfxvU9ZI6NiDcsmGyc4Jyy
lhkmfGUkkrn1xmVRv0afqIru/cFQNtEOPFzqFrj8XDkY9Xe0HbaGTq42yVcISvaD
jmWjWRGzi5qSxrd2qsEhme9SxFKTs9UFQio4A4QmVPZtQf9WaeH9X+UoH5fyNuDG
pW5cxFweVr1pkS0VRdIBiNV71DiU0somchZ7OJPjB1mbacBLUtYA9nPd6E4qW0cI
QaK8zLaDjTBgM+DtsaItoMaTlh6COuO30TW0e+4/u3X6GJ3d2bd+WTGpKW+FLSKw
x3+errKGOlbDeDyS8ntoi1Vyt3tX8BcK2anRijW5lg405wyUO0+X6It6tGUWp8Qe
eazF39SFfw3KA7Lr76Zaq/V1PuJQkFfIMnlZI4+smgy1ckLGdwDmdJBYy7Heb+nH
V5zZ+HUGrGFQKqFsqnp0XJ0Kq/443RK0W1cD6E6VQLo5qPApMtSXVN2yQdfOJUnU
0CaeGemjZIJhGgwe3CGzfjIiXr21QzApygQn2kUBnY2GWjuAdaS5j95m8EWrCEqF
occMhz454Er+i5s8QyahTMp/oK+Qs+BPfnzBQqL/OiQ3w8yCAyldHj77u6qIhdcW
WJKHOnjKx93U8EVMzps/eOvHDXzB/7AfuPxwDz+W8NKGbMVpr/bREfEOg8ULi7ES
98nV0Nf4ceP4laWu53Ec23XontR/SV0rFQ3DUAmADMQx+RwzATFZTXL5JSHxjduB
SwMeyRl+7/dSvnzUGDjDoEllfF5l0C664x/gNexhRvm9pdpbIcBr6jTWUupiot7g
Hm/8v6dRkuPqwFPKny5R7AeVRB732myy9XYK1bch6NZ2BvfujBqJGg6S0fDlo8d9
1MLAYgkviZKqwjZU5foyuyy9a78gCi+MQewB3wsgPqBQiq1/Xkvbw/5YkrBdhPzC
gZNDOYU6AcFsmnMK6gOTAVK29vmaQ/Z0oN+HFrgXCjIuQUKhQzJh1OHcWD1hj193
LztHPYqxuRKuTAF0FfGSSv+rJWzSuW+/O3IWNlsWzbbiWW/mv1ZgjOmRLogYFk7U
U/kSMKUPJn/pnXb+dQBF7H6mnfMy+XADX1EgNBs7het3sR9dC23/KBqQiTNeSJz6
3R7XW8RiRdcAOPdi/l68zrH3x0rxsPWCKGVkdGRZ4Ti5xr71ip4n7o760GMl6Zyh
Afwz6NPNjUP7KzYpKgx8gsxb5nCm0ydMw/tvUGsVxLRxH9JW0aQI5B4dRcXTMEtE
/bPiu939yLpb4aTVSCfuBMVtt5k235erUEnCrCMgSuE3UfxwrdJPDGUnINAdHh29
ub6zfyIGNrPQ9APDITyQE1TPiLC4xq/KcM1cuL9lGCVRTa6Xa4UgDsQmGsZc3Y7O
dD+ukIe7Fuh5SP5cxk7E2Zocj68fwkiLEBUHjxQFMuqpOfgyKokB2h2ZdEYnqtFY
7rodn902mPKx6srX+ELa7nZqhSlu5gAd4r7aMc47Cwp49vyC74ctOle4OJlp+QtS
uwb4Wmj/ZHkgFzeYqruqSxrb1EATooJCLWlvXa7qAaIrF7ut1If+idHY5JwXifRd
89FnO5sfHH9ePSOtmCLjep9HEIYteJZu0L4uU7iytnSPcGooVMY+DWTiNSYMuj33
ISlr5epWR2dwF0qbQGeIQJKR7+dfCFa2ISmlAJTmQUKfitU07JDjXaUml2Vlgi85
9GIZZ6FTNsW5tyvD4ihQc2/hLUwI/QtDUv7JNMvcY2zrZGEyFjy2k01Shdqsey7r
/uZ09QCX30A1Bw//l/iowiEMIeydCkJGvuyx+GXHBdf0T7G/bA5kf7b1kFiiSvU8
N37EmOU6FKa7dQL5+kBkVRZrVm1LE5LRJamBoFuF4kJjaZ3UHr5wcRmD2SH/2xMu
E7MVGhB1OsHhvq3Z9QwYATGMRIn6VEle4KMXX57+0CT76XS/1jvBoXwgVeSQ8DNa
sWLvdaWEeMCOXfNJL6yM6lzxvNV8nbjdrwJzoWGV0WI56cyw/0B7AZ2+IjKdfWqo
q+f+oHA0x0kyYRQImgs0mKKJqPrwV9fAe40nPkicIgsc/s5yExP8U13yNmPJVgYL
Usluma1YCwILsIxFtp7yx/b8pOvslqI1jnWgEgtV9SBkBImzADkcbpdNyIt8TZgu
mF3X4hPUhsxy/euYcfuId4L/G8lWiaa/UpvVBkEsfCk9gGpzqYNLskrY7xf+7UGq
/0ev3z2mZbPhn0r7VR+BUkqnrl26d1Fxt3PesyCeZh7VAi4wnzJ3XXsn0IWxq/SF
wU3WRBsXC3AG/iVyJNxULgJa6sBna3h2hHCd0ows6gxy/Ds01fjhRTjXLh6Y65t7
b8rjHraa6o0ksXASVfs+65C90Qe/eqTxij5ti6L08AgMbuv7oGiKTAhigoq/rJtq
YHSKahWtWFZrVmvQ7lnVixl65Q2hrj/pjXRchLSbaCMJ+j48qI2ecCsfNg16kimv
kn2Hl5s36qxo4IDMVCddz/4n57HsnLtHa7ImUf5wT1bdJvIMvgAed2pFP4MTPgWH
eNNUK/kv1blO3j3rSkdpQT4Ules/UKxZypm7m6i+3dgR1rqf1cpVWjXd71LcznZN
mpol+bsph8l0NepqjG270JS0BwDaHl3A22cQmgWtdlOy0i8+YPAJfLRNYNMgvOJ+
UkHNiSNp4NEV5HDRVhB7C14RIfxtIENXh3oGTDy9wMQV0B2HpVBU/qFovzVEpe0o
FRIIf9xYyTqhMScMef1LjwRzWa+5WM9e68YsnI8J2zY6kxlueR4Ou9U+im5vxfx+
x+hlDle69Z7TA5T5BBP28xRJ2zRopNeGsM4k6BsQ8ivzHYdrTQ7fNoLO3TRAnXHA
uol3frevs5P6e2E8+q3dd6Tc1DN10/1CzQ71TZd02zv4brdzJ2o4b74K+8OKHXiD
dgbVkULRTPilH2FcXQEYCfY45Af+nV+O4gjBXC5PA70mUqp6lWayGD8WGDGGt/Yz
LKvSfr8eeBrh54/ZgDa+bbEbTfU9uuoc65QBkT21bGH9I+/xoKxIMVfWY35/9brI
ilL+wu2F/5hRKYrl8XtMHv8yoFT0wK+pQftbi57CYxFWy2aP2EnCnr1Sf7brDlO7
ZJJllXnx4IrJXowRhAL9YOJIeuetErE249Bty0UpX469BvPx1MfjcQwCaZdHKxwv
NwxA7UIU/vicorShRfN8KYj9DBMzd7cEo0J+OMcRw9gd2RCsD3pzmasLi7agBK2t
jyTP9W/xYeWm20pTttLGhb+7er9VgIcP5qA/Fq93ZVbmHSIpqE66lPNKazYqkEE6
kAqizazpduSsqOF345YqbdezHhZTqurxYuHuO9aBniwJm09+OcsVPsGLJBO/KiI9
QsYGK4lz8XrekkYSCsmhpEY05HLSyzhEO8iduAZC+8PEsvHbHI4nFcBCEJIoaGdR
fNPbqxC64M/9d44PHEpaoxZoDt1Xdo8tr5U5+9dyK2ksHB9Jt/7G7dx8KgrKwWXd
BcZ2v2SzyQ3s7Wym6JtrsjgLlUO/cAljoGIUxU/oixiHBn+3YdCSfGDhgJ1wEK/9
b5DIySeju2ZpOe41eNkt9Cy0sCjpTswOX2aOPUpylgckJMm7goXX0XuaKh7NtBJR
QTmztZG3lBuConHFjAq/Y9bPdm5eWKuLnYomCTSiNAqwrrumrBJFWFsoWJ0tZhdh
GDfgKFS74aNBiF7FBViMWTgwGSQRyCRo3xMjWGIdVvrX6fp3eW44lWXFJaH7u9r7
M5AMgEGA4WfffeXODOXpTFcwDWsWauFUzZD1V4yx6bsuKiA+3CkpWJq+w8MXHqFd
PbUXmmEIGJXku7uWGY1kU/kRnZPhC+tNDKviJfqA9HDh8TjB9aS1rq9opE/qzDwn
f5rJB++nH5ShDN+oWqiWjxdeUjSbzrh0L4kY9UwLY4LlhDFZwkr5IKpksHwV+LgX
PxtR496/YRrEsbnieyKkxQ81Tf7zXqWWDkupwicAnhUYgvOEx33fbjLrc8hCgV53
dKEP3H9rQ1nZE/GhwJKhgQrnLVwWZORvn0/wS0ygtxOXM7xlXVVTHUw2fvO7nil6
/6t8Pj3ukO5SwRo6+f5IDmMfRy60Hw19aOqpvxXXb1vWY1Ynw9sFbrGFYjGO++wH
crJkkLVR8ZjPSdt8SlHA2hMM0/wv0G3zUPcy+//mWmlafAS0FeDu7ZVV6NsGfsKk
1HtYrcFdHmpUbCPC0GAJx4A004fC81mpBzswvbwuFVITuL7LrqEshQmjvliTp+CI
csn09Kt919ixAjzZ2OnI3KmOq1/AQU/v/wAUY/+84mR3/bbj5MbSFNBgn5g0OPZW
7gUpQPHtEmScMRTYWWzVcgwwrARMDdWqDOPKO7UAVfgmFXOkOyxp+Q5OXxq7waJ7
C25OGA2+3pplVIz6RO5KVzQR/2W8eptBsaBJ2Eyiqqt+IRoqlc+yATmqBU5bJEU0
k1MCYx2nkGSnz/UcWFRp4GZepU/agrR17KkfnW/+1DNjQ07L/93viPYz7Hu04Min
7+zSlGbBqTY0YyZApMA9plA2z5LLItq1GE91EmHPkEu4dRoEs+iUtDAdm2lPXD1r
dsd9Atx8ZlzeRTMf9nbjscGpPURp4+BXT16pJps3ZcJl+jeqEu58nDf7kUVVHPvc
eQXP2N8Kv2arlgYzbD64pvkFeWhwG0kMej9A2M1yjl7YKVw8Ej2MAXnM6Ue+hI4Y
yrUuAemFnUNfOlwTOHKlgbfo7joZkvD9cYDteKHLpcwBbIcfG7sla6pjOZJnCWjb
wfnUq8og63i7CX0lMxrqYhqiU3nMYwd9HgbWM1BUvWap3EcjsPdBo76zeKMZjdcb
68ZNfQboYh36go1J/1uPQ+rzrznYAs2qXUBOnpr/OCv2uJaZr9A14FTFpVOZhGcV
d3smHy/zOM1H/qS5umOJPm8q+kOMZkHrslSmhNgT0TjrplilR/kOl8xYAviSCA6+
toMNc+psNbxBjcsIOSLpXzbfNXxR8vE6OFqSErIMw/8A5aFI45jLEUnQYjSFa3Gx
jZIj5P1eDeK07xzSxJnNgcjBBDE2m2PBZD12sYZU5GKraYqvysv+hvZ2YvkoSq3v
bf2IgN5bOiL4nx9+dOH4LyAKzVq8IdPq5V9gAzFWjv1I/iTCrH8Hn/GWqIV4HEkt
Pt6wfYdq8gxZb5LxkyfH3gTvz9IzCEvMPydpxb7MlhM4Be4F0khq27Xy2U8UjO+U
IJWNgOJlwtta7WyPhvHmIDOa4Z+12qi+6iDVxf52vVG3D0R1sN1xVPYtonruQF3e
aHvcOTyGASUyVaWC1f0SxvZ+ZAsjg841C8vWJu14/+WD7gdwSZI+oY5uKfzaf2Oi
2mpxe9lEcYLevkIkLsXbNe2eYc2mDkP9rhvL7TX6mcPlCHemzJj8iR9khIQpWyEX
tOCq2dfCjv/5vzCDGorF6XKTUZt4ZgUo6uEbMjhiWCk=
//pragma protect end_data_block
//pragma protect digest_block
aMwMtoiFI666EU25samLHWWPS1Y=
//pragma protect end_digest_block
//pragma protect end_protected
