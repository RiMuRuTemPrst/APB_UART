/*******************************************************************************
 *    Copyright (C) 2024 by Dolphin Technology
 *    All right reserved.
 *
 *    Copyright Notification
 *    No part may be reproduced except as authorized by written permission.
 *
 *    File Name   : dti_uart_transaction.sv
 *    Company     : Dolphin Technology
 *    Project     : dti uart vip
 *    Author      : Lam Pham Ngoc
 *    Module/Class: dti_uart_transaction
 *    Create Date : Jul 03 2024
 *    Last Update : Jul 03 2024
 *    Description : UART transaction
 ******************************************************************************
  History:

 ******************************************************************************/

class dti_uart_transaction extends uvm_sequence_item;

endclass : dti_uart_transaction