//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
Ak6Fv3vJi/NQTV4466LrtwMpMxVhCbksbu5KeSStqUTQ+nBj0CieT+BGjuAFCIVa
rZq/ZApdCDETIWNfAxTx0lBM86WvYDE9TegTyaLZsv3gmKw6oMuVQdZyKtpyqG/I
X5mzcUzPiIMwqrhpxWucq5cwbNhmE3KybLilVBj3FHos1drWPGThccPLRV/mPvuI
M4a6J0K14hSkwjS6Y8G/wbc9pLlBcAEpSqfbOyc7tegEYPA0jc6SyRikvuT6Ff3P
fG01Igu32n6L7jrDgRk4/6d38Yw4vdnctU/d9fvHsmJIzGJYMqAPzQVpoCDHSAm7
IBxRvP8+M5/WqTnUiSCdvQ==
//pragma protect end_key_block
//pragma protect digest_block
a8sFMIClXqKz+peToprPZBr3ffw=
//pragma protect end_digest_block
//pragma protect data_block
Hm/FI4S1R5zXAje2SvlxJ8SEFgvBd7qDHDYxs2F9Y8FAh4fGKut/3oQtaWbyh5Ip
/U92Odo0tFj4UgO1+AzKptgIS53OPg78q1OW/drhLK/yNzblnF2xTnnj3DMPyNCz
bCjiaufZfJEHID1p3e+RXbLk2NqkIzylrl5E+NbUNX2Qy8sWptdbK7g3TC4hXvwU
Zy4ZEO3fWK3g95xKWoC+PpHph/20GAgoCsF6WkNMmSBwxHXux2CXtNEVz4+p13Gw
QxCOKRjSad/5xTYcEF2F3jBBWgazXzMxPclybEAlCkpFxVhDfy/tVvTb/RJkVxlk
IVGY6k1UWhw9XPVHL7RdAg==
//pragma protect end_data_block
//pragma protect digest_block
4qroG8ZGR3FjSD6Vm+Kuzf6fMuw=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AAp/SBzhLw5kRgiEhYTJjxAcL633OxAYgJAxz1hBGV2sg29wEKp5MopY1VHEOp14
+An94CUwMj5ZLIKesiO9tEj8mUdvWfEFSLpT56xHCDoobsk6SaQwM5lDCQSXABDL
7s9XOeZrJ8zFJQaa5YlKcWZ5WgjjX4MQGXoGJm/GJVo7gE8H0jtOEqD8GcUgNFlp
B7h+F5AM6JMeNcLc8g0nXwxY1c9nYSZdEPypbLjRYgSoGUhTY3DGYv95AL8MoIt5
BQHPuSuXbb/7rJrhkTcmXE4lWWDQ/oxKN98qsSNxP1+u74hWzVSnt6Yfng7Nkgjf
21R7ir8lPCZzpswY2GIHyQ==
//pragma protect end_key_block
//pragma protect digest_block
1fPeLP7ockuZBKNHc9hH6jj8kcM=
//pragma protect end_digest_block
//pragma protect data_block
/Ax0T3TcCHMd4uzX6Ltj79zQ3uVFa3aB3BrbYW8qeyLreJv6w9X/w/fv44nL+z7P
KtVWw2S2Z8gk+m7eh+iy5O4g7EQkxmN6UQGsQnmukCmlgdDKWFJD2xVuZlU/XKNR
Cy8rk6bhZvxzkyn1jOWkQEmXoXmPYchTNbvQa0gTONH6WkPi1IYSguF4O0NLlHFg
8pzHa3zqijJ0pxWB1VGem5aOedJOdb/lvibwzRsoOHnx0juby4TlAjJmQrXZ8ZG7
T+fO4sGaQWXEPi6rC9g3vQBd47PSUs81Bj/LCUBq3Lu6Jpm1ofLkX6plyYyFN4vY
RjqVVdkNyRcG7t93NobYhQ==
//pragma protect end_data_block
//pragma protect digest_block
oa9tHIICPG8RC+L4wILb7l7buMY=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
ATCb8YxxMV5na6QOKjyp37YJQaj+N73mPOQ7vveaIDwQx+EGPx7hT0hX2dVVN9EH
9fjM/IiI6c1E9TUh4owpmFMG6H9BdLWq5a3vnPhDQT1xSIOfZW1OoUL1AFHOBRYv
lpP65nn3s/3hEM47mZI+5rFSDTUCjMwCCt6QkdVG64/UUiFpyvyFSZGTPK8R8ENb
+4IYjr1LBZWghDsqXEY4V0TWJVehpdVot7krkH0S7itVZ712gD49fApTDJEjIiM2
fOvwchIFNM7/Yhq/ruRe0LjQGihdYhvp9XgaRuUK5mG/tJsinvHcaYKO6ES+UfnG
ayfZtgI6xPs9bnSnAFfcow==
//pragma protect end_key_block
//pragma protect digest_block
wMvns37rN4yiiBvO/UKCnElLmTA=
//pragma protect end_digest_block
//pragma protect data_block
JkUz4Hy4IWiwXct9iIYges1DBE/k8QuQYfF4j1qLSH/avAMg9RbGt6rPcpaMUO+r
61hrluMQi7Ij20PAc7YOFIM61CwNzZGdMpEZZMYMu6Hw8gBmDePHo52iF2Ffw3oj
lotPLaNTyEvtrPJnsLu2lADNgrHQ+QUuXmromeW2SbnKFLwcX8JgxYhpWLxjwzQF
QMyYUU7wIU8W6jDT3tIVbI44xUlq5KLRhzMrmOCC5Qjlj5eq/BQ1ApDuKdrOlERs
nbKBolhmOfhUL8pjI9tctQKuGIbhhYntYgdhUEKwlSBLxHvWnLCkSZGK4N6hwUzh
GTm+jBnVTbyWLD/OpknS6g==
//pragma protect end_data_block
//pragma protect digest_block
0pTHb1FdgPzdqQ+cZlO0zV8VXH4=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
Ax5QeSmAIVKxpawqStJHgSwUI1Y6A2yOEga1jvuE2JfcBzaLHIl42ayQs9cb5LJX
puvOHxKQB6VMCGEZoRKQrrJLkvvUUW5cey/YWmfGmIIeAK3CQ98bOlG/TK72NDok
0FhwVIxrpK3eZ3J1L7L5VcgRPlGCodoL4YhkZd5/UYs8XvPbKsgCBvvlcsCk/j6o
UA4Oc3vpjLgTAjHmdcOhFpUolWSVMlLqGhIluK768TDTc7+CLr8/7U04IY4RwjPn
jmqCE8hi6O+21kThvidBDejXozIq1Zr9aS8KrPHQdKwVkZIMo9drpL9iuBOw5YRj
PfSPHAKVRwzGs/HhzRqROw==
//pragma protect end_key_block
//pragma protect digest_block
Oa96QQnAA0F21x5j8zL08WmuuAc=
//pragma protect end_digest_block
//pragma protect data_block
W/suEqTp4Ez80SySl8VGmSQsgDmY1IgCrFwtJgVaMLpcCndQcTETDr8w8k3FE/Gp
gzEWfmYC7rLxV4V1ilO49+BMgqRSojOI2yQFksCAMcs+JVgYyiyplx5TikaHTapM
DBludM0H1V4AOACwnfEt/02sAnNxF23fTZjt7w0Baa418mr9PDOWORYZWyRC1No+
c7bOfKB+dsTvwqNe2iCIh0Yb6jNBtiJj7GonDlnop+K536NPs0MfcwrSn5ELMEA2
mjVrKVtDc9tWWvHF3SNX8M2gG6YpF8TpYQ+TnSmaNxlls5kKDmKB8fvQtrsgoGHJ
kitbZEiQsFP97izoK3H7YGWKigdCDwd1MxEAtLEy9p99RBR/wp/Cj5gj8+VgIbzc
mku6+h7oKxOlGTs2i/+YtGEKfilRXlUoKsiHvM+NQtHxSRzUdgfOjhKKaECb6Qe/
1Av1NCFT4Thr6y0tS8CVOGZV3mH3i5wjZiKLtL5A0/QQgZMMvZeOKfEJ3XGnYfRS
IJWM05NNrsoUFrT01iNK4o1FFoBnlOfLcgb15RdF0kO8IubrHYGDTN9AqSBHvdjl
zjTZwJpfRhzZw8cAlta2USPoIIsGqotTylvUqCFSoL00nCX4pJm2gl0kZ4Vb/nSL
WxEKbLvpx1HGlvsVRtXNXyPofW2NwFxQmV+W8jKapDEccpnzIoXTvZwAmhJDdCPe
WCEdv8TYPfpEcsrmrSvhrFEZdMSfe6DFHHXzekANh5bFtLaE1A0idMpg/JhQMqOf
e3P0HsscdLZll6scO07JyAvAqjFMQgrscMGRkmyLZP1L6iQ7jtDUlqzQtSX3AfpE
cE2IOeHkmRJ22hM8lwH/WRUK2We/e6d1v7wOrxIkQd0FKCGh6C8auhab3C64gxUA
ubUs1aq7ttxwS6pIJ87jJaOhYZMiL8xkF1uniL0ma1p+nEGVBA5n+wIkKeH5ycM2
xbbGi4gniX965MWmn6zUarI/xLXJ6aueq5ISR9KE9XJI6qj63MkS1TzSClRJ5XCz
7QXixiIi07UG8C1A0Rtc64dmXnEoux2EOpPxrOM1EsLQWdM+hsZBY3aFJfDK9Jyl
pJZYVg8WVLWDrAaIt/sISfBEF4KYZXmgt9QYDXSh5pe+kdomM9n+ipwKd8qu418S
6lUjeDXkZOf1+K/66HVfhBHKRM822BZ0bS7xyl8LVx2rGsI4nn9IpmPvl+R5iy27
JX4BuSnV6HHK8ahFni/Kmp/x1Dx71lcTSP9667DVy0qL5XzYx2KAA2t+wg9lJDkH
Cy1+lItZPkdqKeifhF8exzdG8mPlNudn/hQ9K6BrZ+fNvRxcNmioT9eD1iNsUloN
q+g0gaQ7evHVxjAoRUznsmQkII8QeHjA5eFfYwMYiKRl1TSVOylskz2B4vIdjQhm
DkJA18eX6R4t6v+SjdDzzrwLK7jpKX28T5teBHZScnUnkf5/EEcHR5hxXTT1Kd6k
J5dzPsz0fvln6N6rhb3sITxkjSQTb99nUwvlRaxJGWEtE+9XWmdQyZfE+K0GYalN
z+LybULE8v4ifujsKMx1erTPDOZ+IfxSRg97+C5qXEjxDvVT6i9nMUDyzenJpwWf
5MI39B7aNDCtzhN/aSr+1oKKvbMk5GeMQiPU/u0JSXUgMvV9x6Xw09b5CNl3TQAc
Dp67dZ4PFVRLup+RmcUYcYYrfGL7OJeLlI8tneYTD9PlPZO6YIZP3AEbaMaR147P
wKIl220RYAi5+IutBzodpmma+eljtSrRpucoTOGV/1hTJ4fCmrBq6t7GraXVTEkV
z4KYj8YbnGrmuyWNkte0uYC7C1peuGQn2gScL6UQShlfxGS1Gax59DihCDm6fEZU
zDsTve2/XG4e2WMADXAdF8iegEMRnvnPaaDtAdQ63VuYoCpC9iADHkd5GyAxptBe
2y0akQNOsg0EadhzjTodAb1kniM4gZXSwEta9bkE8J8ehz7SdObMo0MoN4aitfup
SW2KC9kOLXmTvpzaXpE2vwctmSO8CUNQaquXLWRQmCZyK5QwPZWhBLTZgk/AaBrx
xWupZCZWCrOOx96ayFrZjmOvUjW7IgCcXAazV9d5ZVt0CTy3wn1tf53GnHF9TMiC
SmIwUDIx2yms5m02h7wq1IElWsUZc2Mq0Ef1dK/sTOG8mE0JsLZJgtwvexeHzZzd
+nlU9E1+lL9yHDfqtply6qQyIIQZsCs7Q3Lv+Ha7c9z438XfH9On1HC28Ma5wq1V
lnGoYJlTnpwRZXXn1iAT8WEZFd9d0Cnvj+1gBgF7k7SjpKVTTC0Ni7WVR3vwpc+H
O+qS/xdI5zPjxd8AubkA6LjsaR+dDa2wmlJCiQLP2+3+BXoD4N34K/ifPJICdHRS
05MNUDp0OClIdymrmCG/0YtsZ/4SZ3fh/iP6ZbVqglZvwS2ZlN2XfNAe2vgkpkmT
DMAhlwiofevA5Flc14sHPuHeEMCrO78ANwIoQP7ulXGVclFNHhwNdnOx2eZInQ1Z
gIg3KfcC0o/qoGB9k787vo1ttQPWw5mPyO3DUb/7497JtRE0RcxOUmaoAMV19mTQ
5iM57ezA9LNiPet81mwsil2OGPBnri6ajCbLfidKJvwrpst11zVpUqOxRBHkfBms
XFlQR2TupvyTleLgVWF8+Qmtm2QOwvvwEQnbGw2z1tQY93bYtO7r70TYdg5DG437
GOyHykAL+q8Ncm7ytMJgfCfNKY2yM+0/rs6au3lRC6RbXhpzcLuXKElkjLjkj0Cj
vwEizbMJ/XGKfd+fIx/j//hNB3RdSYE6lDI3z537avL4xhUpdZnQEPORsvvnZY1y
opYksaH3bX+s8Ej9Ng6/MhYoHc3wy/4uOsNra+52Q7PD0yijXQvn+H8j7665pOWY
2SvLVDK+qpVKoZFgrNO0SNzloosVpMPAJCoqhJM1lQmm5tS43Vl7KarsUHJdMSW5
/70IXcdFPkzRG7AG8sU9/TjA1/u1xM/RpVYRTULowhbfbka7AD/FaTmxbR03WoxZ
zseZaMS7zcpZLJew5tzlKVh1+xuz+zuJHn2FyriiwPmerMmSQTTrkbJiXPvo1UYe
INzgCoHefMtxLhzyFnKb3fK/PzxKAxmJ7QZTjCk/BXh75v4rGsuT/0cV5kB881b1
zewlpJnxQWBKUyCDPv4D+Amu9QU7cNwvGP3CqgpfvdiG4lUHgi6/+ER5ek8VoeSs
6f8adV07NqxnjOjArk/fxC7JVr82Swk7ndZkLW9H2jC0ck69k5GktHYZTTROaoiB
/BWZ7+6Pr74AgfwLkdNO/j3lwBFQCX8ByraGDtt44diaSVcwpxUVzXgi3UsbFtn2
ObkrcC8sPtZW1z/DpI7VQKwTxkw7gL3s8gpURg8nKCkaiMulrtFe1t/rncjpjKEk
6iHpz1GHuUbwizcV7qh2Mjptrkp1v1J4VWjNEqqViklZ0kyoQHTCjzX9TPL2qpq2
HHywsUE0yYJsQtOo81W6i8igjSEQ4/7yHN2fvFyHXgvsn1+3DeOUaDkTDKuCNJVz
3ToRKudWK1Z9zW/eFTKEb2V+ROHg1wLkIfUinDGVbd6TKIgjvOr34VFEbwDoWcnT
w/Cv3qx+78qhVCbpGuZOnvJ5CYaccRyM/pe9wzMmVkoYzm4uLVtni31hVq8NqJPz
kKI8W6fRiey9g0ocW3Rl0whFvdInTrOcfj3tXEdu9omWRSbheM7G5QOLP1x4jJq9
L3Zp4fenLDmdM7544oXZZ3nj499eniEWwDgDEZRhL4DH/e3/jb3+GeAoD3uxZB2w
8+QuRINKNPPlhQI3/N70I5HzgfX6rINBwZoeFIZTkEc5vwd9U4OgN6kLKVleTSQI
MGxReyE35qebcrmbkyKfzQ12A2QM+cOBt4tODPt/QbmQaWkoOMacBC7JG1RNbWmE
6lWgqhgbTaVXs3xEJzD+voBLJOVbdTnqykyi0b5t0og/7BL8SB7XAQ0754qXmMag
tzbAHKLr8xCdHO6/GverRqW3400YC5RK1Io8xYGLvwdH16cTnBsHaEb1LjG8Im0n
xLw895n2q3xI6EzM7Xcc/+axD57pQx8ZSo9D5LHabIz7zXSR6aAErASrB2GhoSap
mxx6OvGl9VXHKSCuYY6gqOxO0TT/m9ajknBvy13Wk0oOyxvDpgCNZQCyoji+7+d8
bNyCU6HsgsqYKCR/bTQkRa4AshzA6LGG1YpbDyefX60z/qYLYA6MIBH/gB8NRuRa
NJrtzA9CTgpTegvgRXrMtGMEbrBGhFjvMstx0k87hh9CC596Mmr9zI0LiUq1KxML
xu+wcPRbN9D1FfNKpBhBWPw/YYmwScmCCV5EAt8CFidEcPySuoOR3Ougpk8A2k58
YkYRnLEac6pIvj/ZzkPmUGHDOPIaP/STio3YyHMT5fc+O6hfv/T+IbQLMgJES/1u
lMS/Po8hx0lKKKAvF3cmXnvCNkbBHCyv9o43pC6bemYQFCeNEsz6w0uGX10V+Jna
37seEAOrrWM6gw2aC+ycof9IsppNQ/M0cGClC9JQqkeEuNkUNFpii+8xG7DoTkKc
hCEgS5Lfq1tYfSWXXrGyReifNKu+rXGmhxY8zRRZt2q2Ec6PvlNjr3cAXTpKTJG3
7K7oyenL3aBvHXUBzwepVmvv7zcaZaeW1ic6P6Gyt+wmCGbjWTMRsoo0aW6eangy
LzX+pouIlT0r6UDG+DtGizjSIBbvzfCwHWrbR2szOTWwLoyY9mRzT0qNrNxnHu5p
4ivb7J3dyBT3EAoixHL/2/K+bCrbPMkoAsoZjklU5u+oO0NFEBM7QNozvj5ptlH7
LDkIfcCECHlKKoXA/E5IRcejjdabBFRCkRAt8oh48N8iuI8uumdYuAYpiNIDqAc3
KhmeLce1mhCAdOXmQq3WTX/x4IzAuSOEP6QJ67G2/zIroBohbE9Bv10yQ7HaG7Xm
WCXTygiU4pjzAirxTsUgp+F27yI5cGjEmNlStTy4/w/hl2TbsM09s7yk5ev/cmu/
zXeS/xd8OD3knun/OzHtB+DriWOFBBOrfKMav87aA9LHdwAAr1hKUDr7leAsiXKT
wvyUqd2Btvs9RvIzWN5qx7G225TJaHp1D8cR6q8q4UpLdRINBZw+DdO/7Zq9Vjvw
TyuA6Oi5UYip0XiNLcwHEzIrChHJGdwZvxF7SRLWxdDth+VVcy7FXx8ZQzOsXhAN
Lt15/yC2W/ARwEam6Rqt33wl7Su17XisSv4Po16yFqeU241MvsnZ+H70h0tS1BQo
4cbQvWqV7wiUCKx3tUnmbGQnTzGqS47JngLN8FN3qu4+5COn8jC1nsbu5H7EE5wF
4mB5GNN6fmsIWRQfQWsoqgTO1do0FQlx7NM8yYXJ52lZ8YD9iSH9M9opd8Gd32xl
IUAQ3JzbvUva1ISpmfhXwIGujLz73CuSdtCjZHdE0oOPfv1eE8bHvLe12YAOelIr
Fi9hpTIXsJmGT9YFbxoGImSgPa8k0RvPEol3RH69EIyw8akhw9qer5RlYbwaqX8m
wtXMRLF3+WUBN6tvvZ+/gpdW8m5vv3QGeH+EFxYyGr5/OJB0xM3thr/GXQjNjnpd
RAVtghAm15NBW7XTdRiopwzXuNlZ8KUmNbT4mg/75XpoQNUg+FQNPjFtYw1+h/oJ
3g6s6vJwCIaX8v8xtAhxOe35VMqWrVhtw1n87pvGNMlCLTaI8ynAh8FWdAP7Fy8i
YLLa4HpHQXcwXaWwei5u2rMvry4gsw0dHyGIb4rWtixFpnDNdHUeY9FHznkf2nPw
1WrE9ARug9CibBGItFGkOjM0Y8ThThJJDo+KVoaqfuMEpmYay0vwRipCsBVk8PQu
XkwnFRXt2oO17Gux8EpLxCU9gjXHCZotDuRET8GCwbpP7eu4krHndp2YdjzfW2Zs
GkyqbnNuQwPFnCUpl5MR2rEmgene6AoyMoyOJ3q19srGmrUcEhto+1xAn1Efhop0
hHmWraczO6i9OT3baRXnmRPYWtWal5GJHzs3Vc7FsBs5HorRzDBoXT+IVglnMtGe
+INifsGBrUcKjNYxmEiHxFtIqQicxJ4bT2YSgPkyQnwFbF87RVK7FPF2lPBGFdr+
TyWAEdqDnTND0gQ3cwkoSt5p75Fi0t7KDhnEG4T6dyjGduRHIOCTQlPuUV8YV4V6
VlTx472NdWok1EjpSx94gRoiXTi36gN+X1RTiyterufykLqfbj35AVTUoQNBwPJL
qzZo0QOkVmzeqUTSy2kZyXIYGvcfWeHQD59eK8XBOZB+H4rZLjzxMbQ1dOC+sYEL
f2Jb3e2ZYOVJ1/HK3ukSN1CiZGzrYCpBsVX8W9b9odqYVAIjlZ+HHYRC18RTDXsQ
SwOzoFWv3tzGZV7UDNTsBKRmiLa6oGm/WDYhaHzKAbs9W2cn8vKDakZel7RgCYUz
tAGxh8s0QcNYMYRCvZY4fuoRD7Pez4NNPivrM2ZQEnFt3ps2vF+oi1tIi1UF8o53
c8t2wuB25MpU8NnlpY3DUN6a4BLmeKS3av/vcRuotuYlHvyKAMkm5nDOrsrcvnFo
3MJXAKAhEhD+nJvvzL3SgBz2VOHh9gBbRXMLPetFr8M77wx/jqOAzEGal/GyKeAv
N1/xACmatTFx46djwKmhTbK9f+oBFkSyeLH7RAapLPJFedZtqcLivkLZSNlKK8dL
pC6xBYCY7l1EOOD8c6Lx00mWeA2l28TEiwgFLLwx9CVYlmqaM3Z/HE4R1g8LXMtO
UDkpgJpYMyL4SP5XxTSoldmkCfRD3acVBy4VWGtTZGZF/DVfZjtQ79iFQZk2ri0Z
KeMI4zn8u7pmOAgVebdp14pXYyaNGnIMhmwlE3X4wvFy199oGA29XMwkicvXefrG
0hf7w9KlEjKWs7Jp1HydkA8zikow/PXgo+mMwHq5F51SWGYUWyMgvG4/G111mWmt
BmMWp7r7NZ7zQwWTlBnJ8VpKP2LqMqErMWd1LkGWLdwowmQnS8kRPnmlwucEDVAc
CBCdmu41A+uqcRAtBXj8/FWh98B7S1e2JQshBNV3PXFNkoweMuTuDewBXB44Wjxm
kzFNyDXOlZv2D8g6eRGrgNMvbMlJMCNcvtrmb6d5Bne+/0fPhqdTevBgnB2hSJja
+UXhx7qk2Wzkf3R8Vv+8RfTvkGIczeOTtIXPH1VQYLp5zbMd0ddWJNdRIkkAHh4H
OXghIZiiFmAAoFXSpDQKGBQdaHGir+hYlVl50G78vG5E270R6M4lXq+32oq0Jrbm
g+xifW++Mv8Un4/rHuSgykTy+Ifh+Beymf8LXUg4eXqWwGcJShbGS2qmclA2EZgF
QVCZ6F60alodvRzoZJtYggUJv8O84fpM27fQ0+rfBLAqf6nVn1HMenMRg14yGpXX
6yrV4IjtlCfnlWOY9EISQL/7rmyC0Pp1orwJwR1UG4qEVDqw5HC3mNR7N9NVRqZL
6Q3UP5N7W4lCKcEirhXXZ1li/G7SFFM5kJlfiZjuE5RpPOY3CmH/0cKbuYvzeMsC
GHs7rI3G9Z3pDQ16SajXZF6cxjiMYYzD0ExYdsqUW9twYjdstCaxj65M38QQ9I29
68yH4KRolthw+JiXvBgjgg7swiwJNAJddvYk4BJ3AU9bHalL2Xn1lmJFqmVM6Pk4
SePahirFpQIJT2Ahw9TS+PmCekTqBQht2aACqXiPcqp3WK86XEERjeG7p6/Z3aO6
Zf4GYEA32pcyniMytNNQg6Me8VYj8prOw0u30QFNuh6xcj9Y7KZWzz4/i+W+5HCD
IfYLaHMua0C3Q+zJvzve6vzWl51HnGMRdBsroa93dVUxEQIIIoJpTESKq5M/xBPz
QnjhlRgfCFb+O+1p1Z0Mf4WWiGyPun6NxID3VHfYYQomC1gbZZx4Y8IEtoazHxsv
AXxNJrEBEIRjo9l9A0jy/pEnltp6THDr5mhVMZucf/LaFBpXrIm9DXIUlcbPLdOv
QHLkUx8ZGE5+P33w33NcnOZ07Zo673vl1JRW46MD5SfXHymAuDZa++zajBV+STkY
E4Ln7Mk01N6j/+KPUN/GPhudCbQOANPnEsx+Em/jXk5hp7dRkjYFSUEM7qaakQAP
Jlt+EIfWlPdP3kkKDio1Xv+ScHLTGAVv3iBBHZf1koTCSjSO99s73spmTFATbZRv
EQZ9J0R55cjpvMFxAT31cdW60btkz/gnXXeUQKV50ZHaPM9qsP9bKRZQP2IYSTvF
RFJsOgE7RzpvWd57P1h5hs0pbK/NbYU0Al5mQd3G6A6fU/Ugww2QO4y0/0bwuXMI
ymMSbxDHYkBHQGV1y/GF/uATWqpUVXTKc5jOOVO0eA6cxIPXVAVZsBsLo4c2EyZh
x0DHqCuUWp64ZWwXTqorNkPRHNgCrXNTvchX1krostsebgVCjkFDcLkVXl5LJ+r6
rMmY5iu5w1uludAWjrjHYJ5sCzYmAgVgtuIoSKRXymv4qSIh85eOu643J/PRqM3k
8XtXoGWzJGELtTJq0Ct8Uf3vUzTNQs3C5U+x1caVCBZYIa9RKm3zwpqYfZ1d+I/A
IvldMXYb3cz6FyJp5lt8z7EKeF8sm1zRjkl677gvy0yXetqvEjfeoJmX26w1zUVC
Iqmp6Loy5nxd9BbQ2m0aIyZqhKsomGJYrwuEAt7YbRB+9Qfmq3bagUDf9SfcBnH2
y2t64vkxxo9xg7kQKXyt2ruxeVeFxLzFmhfMcR13DO52IM1KgxsRuHUs0KcBbLo7
S+IVyBGegSgWq7QpiusiAEz6yRrgZ5or3/kORvYsyW8eT3YS0JRmzjFzN7pMfbjo
DVAhsxDF/oDV1iS1bqHCeXc5iPLBtppuSlRTkpnWK27kk7IGM7+bkK/25L1JQPUU
+ru1eeyX4j7NXM4HuOphTgKHO+uuddHceRosWqdYP1ytxj78TekzSpQKu/u3LTHV
Uny2AQrrRxuq1za4d7K4g6xeO1ysST64lQ22Nw3PJfy/fWu/aTG9o7X6/2vlkLTC
ZCAcjox6VFGj6BJDHSXGsFi3HSaC+6KFP02TyYnf9SkqgG6eXzzHzQioSJK5Zgj3
HVtnQglvsUnlGiwgACYNoxMS6ydg4qgmfzM9NIISB2lRLLdnEbLznfu+46Uk4Bls
QEBIhmokjSC83HYB0nsEqUlXCh2Kq1xSWn9OI5uvcSJ2McDm3xk12Nbt9ErKcp49
f4TDcuyIKub2/dDyIO6VJ4dDT6pno8giQ3JydUMeQ6cYvg6lOMXGCJnt4m/C1gkM
DvECJy5uSJveuYg5GZ1j47CxW0unTEIVg9fjQE3Oy2lxKHZpopqgmbvnfhKtyql4
P2BS1hp6v2aB3MPhKkzfaYbv2cInRIO7AvSJ964CsE02Y6bYB18FuXjR+ASxzhTE
4frdCrFFjI+XKjDbMRVXwJf18OThoJlLHlXVF3NGcAR3ivch+qBfj1bkMarr4IKt
MfV3wWnk+LEzpQSpqip534H/7yCitrOYd3L/HD0ddzGdtnuzwFzTpEemlKBPg1YA
AKHN3/ketIsi4yPzeXZo4gv+A5h0zhjklX5vdYrfXAL9HOojm+69SlRdoOtRizO0
yAn3zBy7ogf7ZOrFVpMneNy5VJVnWgxjz+UOyXPVFA5hyPbncg08J77Z2cLqXNDW
a/T41VMeTzokIfF0YIvXmymr/h4ek5Azvxm1CuwBMUHAQVGGRR5uDYzniYZRATp+
wepRvx8sFATapgx3mplYdRNXjbpiJFqndQVp/jNz5MtaMpqUKLZtxNZOupvAs44W
b7dqbcIhbavFRNNtjr7hmqtZ70XeeAV+qVr4qX2MluzrDTFl+JTZaE0wn9mH1SNs
KPLiIa0Ov7NMzFhYJJBDfYCMekoo2NWeZxNU7OxE94yNJIHETlhvwfm7etAuOHmj
AFKxzYHFpBckAiAS/WI+OGxJUFdtaAyrxA/xG0lS8vURhr5cMim+r2X8J6y0rZn4
vaQdNa8eiFVaCL+9urFVrHThYj9gq1sGuA60G9w91vaXKQDQ7vIdHvM0baudguJ7
1RsL98gBb4VoOIaLJhC8r/Eng3/EI+dZhoAGWQsec4pcB0YhtbYUOL9WCZe+rFfQ
LG0x8ydx1zueEp30FtnbpK7owc14hNx0ratvaUdWagreJieHlR29ESw92FcUWyf2
v4JA9pz1Aqo7TB/MU2eSRXn6gdMpu6+HQwWI36uMNijhdh5HaemvffbEZFABR0Ev
JTzCsDjJMl1QT01JpMjYClLiW6EMSMgRWhxsG6S0N8Mv5pjF96SwPBcN1Ts9aS+1
sMDeVOQZAV5myc4BgXxSowWfIojOe7gUZR8wicQsIxva8ke7USw3/OedIeR6ROQA
dvrMGlTZ31hb7SwSSOQ2JXGaMxLcZrqaPLR+G9LdNBIpKFiVcJAoyy9JImFto6fu
Q+GZfvh8SM+pPzYP+VVRoPvdb9qie49AAbgDzoZxHfFz8d0rKYZElu5p6cCCRqZO
zXBgL9cBUleO6tCzuGp/D9VB7JJy6/30UEXGuUvOWIUhNsoe0GqINZ24EsYHwhiA
8nfMILQQx4RmX6qvHqroR4ZEUhKL4p4giwm/4ZOQVvToEcsjwOoI7wFiGVftvAsX
8LUszi/JnpfuU4Y30umqraaTpuPV4bRVKW9NNPzR+0MR2BfGe9botUntEMbqw0FC
zbfvGddvKjZo5188xcKwjeJCRD4X6j/TJzAYkjwN5JJe1m8AubQ/urNabhNpbE9a
9pHZLqVohP1UalCn5m8VM3OlTO1+5vL/AIX+QKCkzTnraQ85IJA8G5cIfl+DRKu+
yjvLlCIdTV2Ps9UKPW0o752riUZIDuh259wXUUFnUgKLCbUht/8i/mSiYiP5rJMW
9xeLBrqzNz/rGbIDURnFiJ/qcPmcVvMFd+ozIpIeIa01I5LUXXFg6j1sWlT1oSLS
O3c0vxialWFPdoVIIdZaSRvl0fy0jz1smew2y1Cj+03bc8d8UvGgaE4BmsE9oVmC
QNLi4vjZsJy6MpshcDq5Bn81KmdztRbHfqqFfjYt6H5E52vWxtsNHNZDHccJjhD0
bt1+Bd/tbkwFIyKrrz1tG83Q92YvHbWEsK1tslPV4t3itatwgmlXYi94ioajU0Gd
4r+uv0cCfjc4YSZTRNQB0ZgYxW1Jz/8l8jwnS6mlZAWwD9Ptt6mVi2drGbM2pzwd
oCrw92Uogzoiq9O99DgZCDs1OrkCZ/u/pYpLKpJFRPu9BQh7QFymNb6r71MN1rdm
o8mBsTI/bQmRLxVT5WCobhU+53GXHkP9S2a61V4eedJY037ypwpvFDLFLGQXSlvT
5t4lijIz8DuuZ8Ooi5mffqcGZCT3CAsGLZC1udVk9GzlBAqjeJwSidUcrMiS6C/m
iMtd536ZNfulZveTZYDePmZOYDMLvycQOCp5bMbA8LeBNUoUvWOXeasQtHQCgZbn
lJ2b6oBV9Zjwf/dHNB96yhLxDSgO3Y4TLQdkjxZkTtlyv/CtDZWNAkgDDgYlTMVk
XSHaW0fgLMBrQ+fDlEDqoYjJK9PiqvrM/RcSxJhmiZTsSNrXsRABeLGQCjk9iLxg
LF/UJ8VQPVHa5oqV3wYym9w2qMjEudvhlFOuUwLl1R9FxJ4tQISPePuNXsMjRmKZ
ZkML0Ijjh+pZ3P2XAnQHdrons0hXN0iIah8kskpuv7l+YlAgjRAmD7uBixc1a9YW
a69mu6mWUcZYzGDtl3dV6YIWWfOS/15wVtxrMqr+dgLusiZg3KlQ3FmImBm9PD/g
oP0V0ZsDlKCqaEr2WSaf3Ny3ksngWzDLDiRZkM7rUeFicrAS0+IA7wg/x7BW91op
hyVG1UmwcQkMa5tUYKTn3sXcS8Gn6rcPqymaZRgzVlbUknC7ysbpVqGDs5r2H1lx
jOxUax4DJ5Y+EOqCW+wlSGONw+K++VC0zKtU47T6VhcAXJuDJv21dJJrJyAaBeoT
0/mSIpc2kQ9nvm6LVlNDtzFK/jTSmgBelYIJkgEZPqQJVV6nbCdjP/Fg/jV4AoFD
bmL3YyXOOdBfB7JJ824h1xt9D6cLr9EUNn9bfCF9dasUdFrbkdU8mGodxmw0qjG3
31ewpLalEQZXNSEkJsHB+3ZT+eAN/PyoMky9Qaj82qu3x1EGiZDPo/BPSqJT54gJ
THAdNrLxyanR6sVUe8Ur8zha5PvkcZaWE2vCBf8i9IhIbw3rEBmws+ZagCdgRSUa
//pragma protect end_data_block
//pragma protect digest_block
WZ9zyne3QXgTadPyTJy2q3GIxhk=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AGzVsi2gqat3Y7/kdnpG3JRmSHAmEiRNngqFkDay0FtZpuFVXTmor36XzmGrGH8W
g+QP0qr/arHb5GuK1eeC5VkP1akm+W9JdrAICSmqO3/UzST5iT/07+ANVmuz3ABi
pIO3DW4M4toEcXTt+XeQFEt3/QWnTOPILOt/RT2UCBrbTA4CpSjjlaGmJ9ZuLv75
3NmUVnCKSMrtQ4bQSUU/VjWnyGFWOl/XL7fLIthF4S/zr+J8T+/fDCW7B9WP//FT
JLYMsUNiJAavqsuovxkyU+7rcURWDg6wDN64frMbs8lB4clG0k/CLCrW7292KmmR
HNl9VXibH0FN0z17F8Rg8A==
//pragma protect end_key_block
//pragma protect digest_block
kW335nXE7P1QDuV9E602nSpH3vw=
//pragma protect end_digest_block
//pragma protect data_block
H4z3R9ImxuVEvqrGP6vsrm6Y+xl01G4PJqmwKKt21oJRviBzr3/ooG1y/YUln5TQ
r2W09sBSSWQ7SBAJvR6qPlvkrmyFaIV09jg/H4xqTGHdN6QW4JhrDXBvqH5cvnWo
YhpbAnidC1R/ym/v29+zP6nE0yjPgl2jcBl3xH9qThd9FFazgXvbv0ndEImF76YW
YGL8iCOP+asLORkRbOId0385Z8TP1zTZW/uG3HrGYQdu6sZ3hoCJOWTvNnyWnKdy
QwcD/hF/PU9kPv2nC3UA8jkILYSvy9iMYD3roP2yi5CgQAPnHP/mMb+/hr+3e2Kc
zn1jfrIwDKhNKl5nWrAU6w==
//pragma protect end_data_block
//pragma protect digest_block
kwrgcaPWgtHFat604dLxP7xRxpM=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AwxcPhdhV4xtuujWdNKKGpMYxJFtfP0P0/M5a/Y0mPiiY3ImqsnrrLKrmbeNvXoH
2ki6vTFX3iMPmBXOzasKeXVgANJcO1EDSSwbzV/Q77JZjBg/+oHSoAMXe7dRD/uc
sq2lU2Ecju6gX7S/G3iOm+vv4IuYerlsbu2+G0n1DYGrLjhv6p32tJC0uYjHX+Fb
wzWNTnxkV0aSoqwkxFAyoRExr2YDRBJLKeHEpndD1D3oM5GpuBk9QoYJQ5Lf1/6+
HS82O8W9TK5Idrfof5GtDtibfcd/NC7c12lOEIkKlMzk0mR389ba5k/jnUPIN6YV
PFC1tT/y+uVpTQ2i3npCkQ==
//pragma protect end_key_block
//pragma protect digest_block
1GpsSP+YvXhv8iI8Zy8cqsAx0Mg=
//pragma protect end_digest_block
//pragma protect data_block
+KHmFl1I29nDek3Pnew/fZhzkpmUsvKDKnV1Dhqk2z2yi3lBe0CIMsMt5dqdzuoj
DEM8b0SEG4Lk1NKvN2A5QVEVVuxAjXtMPMtlsRbLbOfNNKMyjQF78g1HQ68h1Lpw
VCgQSMbi1UOtes9Vz06NTb9MwDAiYXe/LbeFyQurf1t4z8mgtQHuy+ryvKMBVxpL
Cj+LXzj7Ho/bmAb50JGzSvd11oF46ndhtOrTF733NIvA1T6lmj0DC4w05QjS8iMK
GHVAPHKYgoYa6jH1kFnM+wUr8Bepbhi1ltA12JUT5qQkPYZvjT/Agnk6RXZTY+bQ
ITqr7HOjrlKAwV7741c1mA==
//pragma protect end_data_block
//pragma protect digest_block
nCQfqnVFkDssImUbRg18IQXgsYA=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_2)
//pragma protect key_method=RSA
//pragma protect key_block
AsKyccDi+pIS53g1Dzn8dn6rT468lFMsPK358o94BZZTRSDKZ8pghLpCtHRnu6Qf
tG53T79GUzVhO6+0CffjXqIt/wsYzap9OwUKxcuK1T/LAC0bdakA3JIhHLU9IXzF
IHUWcHo0ZFHMs869ydiZ/GCK3meSasPdOayCawnL4RMJdd+nv23KMEOH4OsS6bWA
3CsjFh4aAncM3BYuY/aPBVzD0P/x2XFSaPWSDK9DNpBbMdjh/PegwYkTduSExN5b
PWucjsD51LaynsDZnWSYnS+kPgCbV2xWTLkvwoXCDd3bQhwr3F41WUVUsDp4KBKA
86aNZYnw9piL4oHhWLNYAg==
//pragma protect end_key_block
//pragma protect digest_block
gXAQnUIxdqHgmIQEd6YQctVW/Sw=
//pragma protect end_digest_block
//pragma protect data_block
23Fm0M9Zv1IHOKEOq0aKVrIhF8a9kOYyJ2dlKoZgMx+UQtmD/F2IeoB4HEW14qsg
/BUmD7D5oD33ejMpuuI2ht+56eRwiaukKKFy2DdVcx81akA5X0+Sin7GItLp5v3Y
y+V0UkSLomXn6h0cbPXvUz7Zz+OO++sCwp7RuO2RApXeFVGFaX1QxHYytwCJwmt5
i26y8lK0ZSgo6DlmWg36x8sZ7Dt9SpnSAWuNn9aIwJ6v1jSAL700wm3lEPPCtgao
9frTRXmnmjiIIyg1WAgnzBP9yudv1nURTfCGqEZJMFv64zJFwBpChj62Xhzm+a/t
RbkYttpjJGOnc3D/6xbUUQ==
//pragma protect end_data_block
//pragma protect digest_block
rO+GNuC7cSJTcK8NJOHxxa9OxPw=
//pragma protect end_digest_block
//pragma protect end_protected
